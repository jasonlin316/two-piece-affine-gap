# Confidential Information of ARM, Inc.
# Use subject to ARM license.
# Copyright (c) 2020 ARM, Inc.

# ACI Version r11p2

# Reifier 3.1.1

VERSION 5.6 ;

BUSBITCHARS "[]" ;

#name: High Density Single Port SRAM RVT-HVT-RVT Compiler|CLN40G 40nm Process, 256 Rows Per Bank, 0.299um^2 Bit Cell
#version: r11p2
#comment: 
#configuration:  -instname "sram_sp_hde" -words 2048 -bits 80 -frequency 1 -mux 8 -pipeline off -write_mask off -wp_size 1 -write_thru on -top_layer "m5-m9" -power_type otc -redundancy off -rcols 2 -rrows 4 -bmux on -ser none -power_gating off -retention on -ema on -atf off -cust_comment "" -bus_notation on -left_bus_delim "[" -right_bus_delim "]" -pwr_gnd_rename "vddpe:VDDPE,vddce:VDDCE,vsse:VSSE" -prefix "" -name_case upper -rows_p_bl 256 -check_instname on -diodes on -drive 6 -dnw off -corners tt_0p90v_0p90v_25c,ss_0p81v_0p81v_m40c,ss_0p81v_0p81v_125c,ffg_0p99v_0p99v_125c,ff_0p99v_0p99v_m40c,ff_0p99v_0p99v_125c
SITE sram_sp_hde
  CLASS  CORE ;
  SIZE 572.31 BY 145.84 ;
  END sram_sp_hde

MACRO sram_sp_hde
  FOREIGN sram_sp_hde 0 0 ;
  SYMMETRY X Y R90 ;
  SITE sram_sp_hde ;
  SIZE 572.31 BY 145.84 ;
  CLASS BLOCK ;
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 297.66 0.0 297.8 0.07 ;
      LAYER M4 ;
      RECT 297.66 0.0 297.8 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[41]
  PIN TA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 297.34 0.0 297.48 0.07 ;
      LAYER M1 ;
      RECT 297.34 0.0 297.48 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[8]
  PIN TD[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 298.08 0.0 298.22 0.07 ;
      LAYER M4 ;
      RECT 298.08 0.0 298.22 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[41]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 297.09 0.0 297.23 0.07 ;
      LAYER M1 ;
      RECT 297.09 0.0 297.23 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[41]
  PIN DY[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 298.29 0.0 298.43 0.07 ;
      LAYER M2 ;
      RECT 298.29 0.0 298.43 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[41]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 294.205 0.0 294.345 0.07 ;
      LAYER M1 ;
      RECT 294.205 0.0 294.345 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[8]
  PIN AY[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 298.61 0.0 298.75 0.07 ;
      LAYER M2 ;
      RECT 298.61 0.0 298.75 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[8]
  PIN TQ[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 292.99 0.0 293.13 0.07 ;
      LAYER M3 ;
      RECT 292.99 0.0 293.13 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[40]
  PIN TQ[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 299.63 0.0 299.77 0.07 ;
      LAYER M4 ;
      RECT 299.63 0.0 299.77 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[41]
  PIN AY[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 292.005 0.0 292.145 0.07 ;
      LAYER M1 ;
      RECT 292.005 0.0 292.145 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[9]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 300.825 0.0 300.965 0.07 ;
      LAYER M2 ;
      RECT 300.825 0.0 300.965 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[7]
  PIN DY[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 291.65 0.0 291.79 0.07 ;
      LAYER M1 ;
      RECT 291.65 0.0 291.79 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[40]
  PIN TA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 303.48 0.0 303.62 0.07 ;
      LAYER M2 ;
      RECT 303.48 0.0 303.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[7]
  PIN TD[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 291.44 0.0 291.58 0.07 ;
      LAYER M3 ;
      RECT 291.44 0.0 291.58 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[40]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 303.73 0.0 303.87 0.07 ;
      LAYER M2 ;
      RECT 303.73 0.0 303.87 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[42]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 291.02 0.0 291.16 0.07 ;
      LAYER M3 ;
      RECT 291.02 0.0 291.16 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[40]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 304.3 0.0 304.44 0.07 ;
      LAYER M4 ;
      RECT 304.3 0.0 304.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[42]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 290.81 0.0 290.95 0.07 ;
      LAYER M1 ;
      RECT 290.81 0.0 290.95 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END CLK
  PIN TD[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 304.72 0.0 304.86 0.07 ;
      LAYER M4 ;
      RECT 304.72 0.0 304.86 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[42]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 290.45 0.0 290.59 0.07 ;
      LAYER M1 ;
      RECT 290.45 0.0 290.59 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[40]
  PIN DY[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 304.93 0.0 305.07 0.07 ;
      LAYER M2 ;
      RECT 304.93 0.0 305.07 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[42]
  PIN TA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 286.295 0.0 286.435 0.07 ;
      LAYER M1 ;
      RECT 286.295 0.0 286.435 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[9]
  PIN TQ[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 306.27 0.0 306.41 0.07 ;
      LAYER M4 ;
      RECT 306.27 0.0 306.41 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[42]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 286.045 0.0 286.185 0.07 ;
      LAYER M1 ;
      RECT 286.045 0.0 286.185 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[9]
  PIN AY[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 306.535 0.0 306.675 0.07 ;
      LAYER M2 ;
      RECT 306.535 0.0 306.675 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[7]
  PIN RET1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 285.685 0.0 285.825 0.07 ;
      LAYER M1 ;
      RECT 285.685 0.0 285.825 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END RET1N
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 307.3 0.0 307.44 0.07 ;
      LAYER M2 ;
      RECT 307.3 0.0 307.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[6]
  PIN AY[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 283.27 0.0 283.41 0.07 ;
      LAYER M1 ;
      RECT 283.27 0.0 283.41 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[10]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 310.37 0.0 310.51 0.07 ;
      LAYER M2 ;
      RECT 310.37 0.0 310.51 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[43]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 282.215 0.0 282.355 0.07 ;
      LAYER M1 ;
      RECT 282.215 0.0 282.355 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[39]
  PIN TA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 310.785 0.0 310.925 0.07 ;
      LAYER M2 ;
      RECT 310.785 0.0 310.925 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[6]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 281.15 0.0 281.29 0.07 ;
      LAYER M3 ;
      RECT 281.15 0.0 281.29 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[39]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 310.94 0.0 311.08 0.07 ;
      LAYER M4 ;
      RECT 310.94 0.0 311.08 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[43]
  PIN DY[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 280.98 0.0 281.12 0.07 ;
      LAYER M1 ;
      RECT 280.98 0.0 281.12 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[39]
  PIN TD[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 311.36 0.0 311.5 0.07 ;
      LAYER M4 ;
      RECT 311.36 0.0 311.5 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[43]
  PIN TD[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 280.73 0.0 280.87 0.07 ;
      LAYER M3 ;
      RECT 280.73 0.0 280.87 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[39]
  PIN DY[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 311.57 0.0 311.71 0.07 ;
      LAYER M2 ;
      RECT 311.57 0.0 311.71 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[43]
  PIN TQ[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 279.18 0.0 279.32 0.07 ;
      LAYER M3 ;
      RECT 279.18 0.0 279.32 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[39]
  PIN TQ[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 312.91 0.0 313.05 0.07 ;
      LAYER M4 ;
      RECT 312.91 0.0 313.05 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[43]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 278.93 0.0 279.07 0.07 ;
      LAYER M1 ;
      RECT 278.93 0.0 279.07 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[10]
  PIN AY[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 313.195 0.0 313.335 0.07 ;
      LAYER M2 ;
      RECT 313.195 0.0 313.335 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[6]
  PIN TA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 278.235 0.0 278.375 0.07 ;
      LAYER M1 ;
      RECT 278.235 0.0 278.375 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[10]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 314.105 0.0 314.245 0.07 ;
      LAYER M2 ;
      RECT 314.105 0.0 314.245 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[5]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 275.445 0.0 275.585 0.07 ;
      LAYER M1 ;
      RECT 275.445 0.0 275.585 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[38]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 317.01 0.0 317.15 0.07 ;
      LAYER M2 ;
      RECT 317.01 0.0 317.15 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[44]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 274.51 0.0 274.65 0.07 ;
      LAYER M3 ;
      RECT 274.51 0.0 274.65 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[38]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 317.58 0.0 317.72 0.07 ;
      LAYER M4 ;
      RECT 317.58 0.0 317.72 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[44]
  PIN DY[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 274.3 0.0 274.44 0.07 ;
      LAYER M1 ;
      RECT 274.3 0.0 274.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[38]
  PIN TD[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 318.0 0.0 318.14 0.07 ;
      LAYER M4 ;
      RECT 318.0 0.0 318.14 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[44]
  PIN TD[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 274.09 0.0 274.23 0.07 ;
      LAYER M3 ;
      RECT 274.09 0.0 274.23 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[38]
  PIN DY[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 318.21 0.0 318.35 0.07 ;
      LAYER M2 ;
      RECT 318.21 0.0 318.35 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[44]
  PIN TQ[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 272.54 0.0 272.68 0.07 ;
      LAYER M3 ;
      RECT 272.54 0.0 272.68 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[38]
  PIN TA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 319.24 0.0 319.38 0.07 ;
      LAYER M2 ;
      RECT 319.24 0.0 319.38 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[5]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 268.805 0.0 268.945 0.07 ;
      LAYER M1 ;
      RECT 268.805 0.0 268.945 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[37]
  PIN TQ[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 319.55 0.0 319.69 0.07 ;
      LAYER M4 ;
      RECT 319.55 0.0 319.69 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[44]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 267.87 0.0 268.01 0.07 ;
      LAYER M3 ;
      RECT 267.87 0.0 268.01 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[37]
  PIN AY[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 320.08 0.0 320.22 0.07 ;
      LAYER M2 ;
      RECT 320.08 0.0 320.22 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[5]
  PIN DY[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 267.66 0.0 267.8 0.07 ;
      LAYER M1 ;
      RECT 267.66 0.0 267.8 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[37]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 321.85 0.0 321.99 0.07 ;
      LAYER M2 ;
      RECT 321.85 0.0 321.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END CEN
  PIN TD[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 267.45 0.0 267.59 0.07 ;
      LAYER M3 ;
      RECT 267.45 0.0 267.59 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[37]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 323.65 0.0 323.79 0.07 ;
      LAYER M2 ;
      RECT 323.65 0.0 323.79 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[45]
  PIN BEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 266.14 0.0 266.28 0.07 ;
      LAYER M1 ;
      RECT 266.14 0.0 266.28 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END BEN
  PIN TCEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 324.18 0.0 324.32 0.07 ;
      LAYER M2 ;
      RECT 324.18 0.0 324.32 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TCEN
  PIN TQ[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.9 0.0 266.04 0.07 ;
      LAYER M3 ;
      RECT 265.9 0.0 266.04 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[37]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 324.22 0.0 324.36 0.07 ;
      LAYER M4 ;
      RECT 324.22 0.0 324.36 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[45]
  PIN TEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 263.88 0.0 264.02 0.07 ;
      LAYER M1 ;
      RECT 263.88 0.0 264.02 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TEN
  PIN TD[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 324.64 0.0 324.78 0.07 ;
      LAYER M4 ;
      RECT 324.64 0.0 324.78 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[45]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 262.165 0.0 262.305 0.07 ;
      LAYER M1 ;
      RECT 262.165 0.0 262.305 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[36]
  PIN DY[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 324.85 0.0 324.99 0.07 ;
      LAYER M2 ;
      RECT 324.85 0.0 324.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[45]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 261.23 0.0 261.37 0.07 ;
      LAYER M3 ;
      RECT 261.23 0.0 261.37 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[36]
  PIN TQ[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 326.19 0.0 326.33 0.07 ;
      LAYER M4 ;
      RECT 326.19 0.0 326.33 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[45]
  PIN DY[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 261.02 0.0 261.16 0.07 ;
      LAYER M1 ;
      RECT 261.02 0.0 261.16 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[36]
  PIN CENY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 327.325 0.0 327.465 0.07 ;
      LAYER M2 ;
      RECT 327.325 0.0 327.465 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END CENY
  PIN TD[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 260.81 0.0 260.95 0.07 ;
      LAYER M3 ;
      RECT 260.81 0.0 260.95 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[36]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 330.29 0.0 330.43 0.07 ;
      LAYER M2 ;
      RECT 330.29 0.0 330.43 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[46]
  PIN EMAS
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 259.54 0.0 259.68 0.07 ;
      LAYER M1 ;
      RECT 259.54 0.0 259.68 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAS
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 330.86 0.0 331.0 0.07 ;
      LAYER M4 ;
      RECT 330.86 0.0 331.0 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[46]
  PIN TQ[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 259.26 0.0 259.4 0.07 ;
      LAYER M3 ;
      RECT 259.26 0.0 259.4 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[36]
  PIN TD[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 331.28 0.0 331.42 0.07 ;
      LAYER M4 ;
      RECT 331.28 0.0 331.42 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[46]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 255.525 0.0 255.665 0.07 ;
      LAYER M1 ;
      RECT 255.525 0.0 255.665 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[35]
  PIN DY[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 331.49 0.0 331.63 0.07 ;
      LAYER M2 ;
      RECT 331.49 0.0 331.63 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[46]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 254.59 0.0 254.73 0.07 ;
      LAYER M3 ;
      RECT 254.59 0.0 254.73 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[35]
  PIN TQ[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 332.83 0.0 332.97 0.07 ;
      LAYER M4 ;
      RECT 332.83 0.0 332.97 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[46]
  PIN TD[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 254.17 0.0 254.31 0.07 ;
      LAYER M3 ;
      RECT 254.17 0.0 254.31 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[35]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 336.93 0.0 337.07 0.07 ;
      LAYER M2 ;
      RECT 336.93 0.0 337.07 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[47]
  PIN DY[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 253.96 0.0 254.1 0.07 ;
      LAYER M1 ;
      RECT 253.96 0.0 254.1 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[35]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 337.5 0.0 337.64 0.07 ;
      LAYER M4 ;
      RECT 337.5 0.0 337.64 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[47]
  PIN TQ[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 252.62 0.0 252.76 0.07 ;
      LAYER M3 ;
      RECT 252.62 0.0 252.76 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[35]
  PIN TD[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 337.92 0.0 338.06 0.07 ;
      LAYER M4 ;
      RECT 337.92 0.0 338.06 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[47]
  PIN EMAW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 251.79 0.0 251.93 0.07 ;
      LAYER M1 ;
      RECT 251.79 0.0 251.93 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAW[0]
  PIN DY[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 338.13 0.0 338.27 0.07 ;
      LAYER M2 ;
      RECT 338.13 0.0 338.27 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[47]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 248.52 0.0 248.66 0.07 ;
      LAYER M1 ;
      RECT 248.52 0.0 248.66 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[34]
  PIN TQ[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 339.47 0.0 339.61 0.07 ;
      LAYER M4 ;
      RECT 339.47 0.0 339.61 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[47]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 247.95 0.0 248.09 0.07 ;
      LAYER M3 ;
      RECT 247.95 0.0 248.09 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[34]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 343.57 0.0 343.71 0.07 ;
      LAYER M2 ;
      RECT 343.57 0.0 343.71 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[48]
  PIN TD[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 247.53 0.0 247.67 0.07 ;
      LAYER M3 ;
      RECT 247.53 0.0 247.67 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[34]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 344.14 0.0 344.28 0.07 ;
      LAYER M4 ;
      RECT 344.14 0.0 344.28 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[48]
  PIN DY[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 247.32 0.0 247.46 0.07 ;
      LAYER M1 ;
      RECT 247.32 0.0 247.46 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[34]
  PIN TD[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 344.56 0.0 344.7 0.07 ;
      LAYER M4 ;
      RECT 344.56 0.0 344.7 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[48]
  PIN TQ[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 245.98 0.0 246.12 0.07 ;
      LAYER M3 ;
      RECT 245.98 0.0 246.12 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[34]
  PIN DY[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 344.77 0.0 344.91 0.07 ;
      LAYER M2 ;
      RECT 344.77 0.0 344.91 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[48]
  PIN EMAW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 243.465 0.0 243.605 0.07 ;
      LAYER M1 ;
      RECT 243.465 0.0 243.605 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAW[1]
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 345.125 0.0 345.265 0.07 ;
      LAYER M2 ;
      RECT 345.125 0.0 345.265 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END WEN
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 241.88 0.0 242.02 0.07 ;
      LAYER M1 ;
      RECT 241.88 0.0 242.02 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[33]
  PIN TWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 345.795 0.0 345.935 0.07 ;
      LAYER M2 ;
      RECT 345.795 0.0 345.935 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TWEN
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 241.31 0.0 241.45 0.07 ;
      LAYER M3 ;
      RECT 241.31 0.0 241.45 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[33]
  PIN TQ[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 346.11 0.0 346.25 0.07 ;
      LAYER M4 ;
      RECT 346.11 0.0 346.25 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[48]
  PIN TD[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 240.89 0.0 241.03 0.07 ;
      LAYER M3 ;
      RECT 240.89 0.0 241.03 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[33]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 350.21 0.0 350.35 0.07 ;
      LAYER M2 ;
      RECT 350.21 0.0 350.35 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[49]
  PIN DY[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 240.68 0.0 240.82 0.07 ;
      LAYER M1 ;
      RECT 240.68 0.0 240.82 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[33]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 350.78 0.0 350.92 0.07 ;
      LAYER M4 ;
      RECT 350.78 0.0 350.92 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[49]
  PIN EMA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 239.65 0.0 239.79 0.07 ;
      LAYER M1 ;
      RECT 239.65 0.0 239.79 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END EMA[0]
  PIN TD[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 351.2 0.0 351.34 0.07 ;
      LAYER M4 ;
      RECT 351.2 0.0 351.34 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[49]
  PIN TQ[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 239.34 0.0 239.48 0.07 ;
      LAYER M3 ;
      RECT 239.34 0.0 239.48 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[33]
  PIN DY[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 351.41 0.0 351.55 0.07 ;
      LAYER M2 ;
      RECT 351.41 0.0 351.55 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[49]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 235.24 0.0 235.38 0.07 ;
      LAYER M1 ;
      RECT 235.24 0.0 235.38 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[32]
  PIN WENY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 351.765 0.0 351.905 0.07 ;
      LAYER M2 ;
      RECT 351.765 0.0 351.905 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END WENY
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 234.67 0.0 234.81 0.07 ;
      LAYER M3 ;
      RECT 234.67 0.0 234.81 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[32]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 352.435 0.0 352.575 0.07 ;
      LAYER M2 ;
      RECT 352.435 0.0 352.575 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[4]
  PIN TD[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 234.25 0.0 234.39 0.07 ;
      LAYER M3 ;
      RECT 234.25 0.0 234.39 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[32]
  PIN TQ[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 352.75 0.0 352.89 0.07 ;
      LAYER M4 ;
      RECT 352.75 0.0 352.89 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[49]
  PIN DY[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 234.04 0.0 234.18 0.07 ;
      LAYER M1 ;
      RECT 234.04 0.0 234.18 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[32]
  PIN TA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 352.955 0.0 353.095 0.07 ;
      LAYER M2 ;
      RECT 352.955 0.0 353.095 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[4]
  PIN TQ[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 232.7 0.0 232.84 0.07 ;
      LAYER M3 ;
      RECT 232.7 0.0 232.84 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[32]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 356.85 0.0 356.99 0.07 ;
      LAYER M2 ;
      RECT 356.85 0.0 356.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[50]
  PIN EMA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 230.435 0.0 230.575 0.07 ;
      LAYER M1 ;
      RECT 230.435 0.0 230.575 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END EMA[1]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 357.42 0.0 357.56 0.07 ;
      LAYER M4 ;
      RECT 357.42 0.0 357.56 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[50]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 228.6 0.0 228.74 0.07 ;
      LAYER M1 ;
      RECT 228.6 0.0 228.74 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[31]
  PIN TD[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 357.84 0.0 357.98 0.07 ;
      LAYER M4 ;
      RECT 357.84 0.0 357.98 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[50]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 228.03 0.0 228.17 0.07 ;
      LAYER M3 ;
      RECT 228.03 0.0 228.17 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[31]
  PIN DY[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 358.05 0.0 358.19 0.07 ;
      LAYER M2 ;
      RECT 358.05 0.0 358.19 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[50]
  PIN TD[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 227.61 0.0 227.75 0.07 ;
      LAYER M3 ;
      RECT 227.61 0.0 227.75 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[31]
  PIN AY[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 358.37 0.0 358.51 0.07 ;
      LAYER M2 ;
      RECT 358.37 0.0 358.51 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[4]
  PIN DY[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 227.4 0.0 227.54 0.07 ;
      LAYER M1 ;
      RECT 227.4 0.0 227.54 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[31]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 359.075 0.0 359.215 0.07 ;
      LAYER M2 ;
      RECT 359.075 0.0 359.215 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[3]
  PIN TQ[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 226.06 0.0 226.2 0.07 ;
      LAYER M3 ;
      RECT 226.06 0.0 226.2 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[31]
  PIN TQ[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 359.39 0.0 359.53 0.07 ;
      LAYER M4 ;
      RECT 359.39 0.0 359.53 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[50]
  PIN EMA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 224.995 0.0 225.135 0.07 ;
      LAYER M1 ;
      RECT 224.995 0.0 225.135 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END EMA[2]
  PIN TA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 362.395 0.0 362.535 0.07 ;
      LAYER M2 ;
      RECT 362.395 0.0 362.535 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[3]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 221.96 0.0 222.1 0.07 ;
      LAYER M1 ;
      RECT 221.96 0.0 222.1 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[30]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 363.49 0.0 363.63 0.07 ;
      LAYER M2 ;
      RECT 363.49 0.0 363.63 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[51]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 221.39 0.0 221.53 0.07 ;
      LAYER M3 ;
      RECT 221.39 0.0 221.53 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[30]
  PIN AY[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 363.905 0.0 364.045 0.07 ;
      LAYER M2 ;
      RECT 363.905 0.0 364.045 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[3]
  PIN TD[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 220.97 0.0 221.11 0.07 ;
      LAYER M3 ;
      RECT 220.97 0.0 221.11 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[30]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 364.06 0.0 364.2 0.07 ;
      LAYER M4 ;
      RECT 364.06 0.0 364.2 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[51]
  PIN DY[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 220.76 0.0 220.9 0.07 ;
      LAYER M1 ;
      RECT 220.76 0.0 220.9 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[30]
  PIN TD[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 364.48 0.0 364.62 0.07 ;
      LAYER M4 ;
      RECT 364.48 0.0 364.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[51]
  PIN STOV
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 219.63 0.0 219.77 0.07 ;
      LAYER M1 ;
      RECT 219.63 0.0 219.77 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END STOV
  PIN DY[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 364.69 0.0 364.83 0.07 ;
      LAYER M2 ;
      RECT 364.69 0.0 364.83 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[51]
  PIN TQ[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 219.42 0.0 219.56 0.07 ;
      LAYER M3 ;
      RECT 219.42 0.0 219.56 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[30]
  PIN TQ[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 366.03 0.0 366.17 0.07 ;
      LAYER M4 ;
      RECT 366.03 0.0 366.17 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[51]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 215.32 0.0 215.46 0.07 ;
      LAYER M1 ;
      RECT 215.32 0.0 215.46 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[29]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 370.13 0.0 370.27 0.07 ;
      LAYER M2 ;
      RECT 370.13 0.0 370.27 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[52]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 214.75 0.0 214.89 0.07 ;
      LAYER M3 ;
      RECT 214.75 0.0 214.89 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[29]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 370.7 0.0 370.84 0.07 ;
      LAYER M4 ;
      RECT 370.7 0.0 370.84 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[52]
  PIN TD[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 214.33 0.0 214.47 0.07 ;
      LAYER M3 ;
      RECT 214.33 0.0 214.47 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[29]
  PIN TD[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 371.12 0.0 371.26 0.07 ;
      LAYER M4 ;
      RECT 371.12 0.0 371.26 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[52]
  PIN DY[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 214.12 0.0 214.26 0.07 ;
      LAYER M1 ;
      RECT 214.12 0.0 214.26 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[29]
  PIN DY[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 371.33 0.0 371.47 0.07 ;
      LAYER M2 ;
      RECT 371.33 0.0 371.47 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[52]
  PIN TQ[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 212.78 0.0 212.92 0.07 ;
      LAYER M3 ;
      RECT 212.78 0.0 212.92 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[29]
  PIN TQ[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 372.67 0.0 372.81 0.07 ;
      LAYER M4 ;
      RECT 372.67 0.0 372.81 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[52]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 208.68 0.0 208.82 0.07 ;
      LAYER M1 ;
      RECT 208.68 0.0 208.82 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[28]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 376.77 0.0 376.91 0.07 ;
      LAYER M2 ;
      RECT 376.77 0.0 376.91 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[53]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 208.11 0.0 208.25 0.07 ;
      LAYER M3 ;
      RECT 208.11 0.0 208.25 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[28]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 377.34 0.0 377.48 0.07 ;
      LAYER M4 ;
      RECT 377.34 0.0 377.48 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[53]
  PIN TD[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 207.69 0.0 207.83 0.07 ;
      LAYER M3 ;
      RECT 207.69 0.0 207.83 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[28]
  PIN TD[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 377.76 0.0 377.9 0.07 ;
      LAYER M4 ;
      RECT 377.76 0.0 377.9 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[53]
  PIN DY[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 207.48 0.0 207.62 0.07 ;
      LAYER M1 ;
      RECT 207.48 0.0 207.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[28]
  PIN DY[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 377.97 0.0 378.11 0.07 ;
      LAYER M2 ;
      RECT 377.97 0.0 378.11 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[53]
  PIN TQ[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 206.14 0.0 206.28 0.07 ;
      LAYER M3 ;
      RECT 206.14 0.0 206.28 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[28]
  PIN TQ[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 379.31 0.0 379.45 0.07 ;
      LAYER M4 ;
      RECT 379.31 0.0 379.45 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[53]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 202.04 0.0 202.18 0.07 ;
      LAYER M1 ;
      RECT 202.04 0.0 202.18 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[27]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 379.53 0.0 379.67 0.07 ;
      LAYER M2 ;
      RECT 379.53 0.0 379.67 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[2]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 201.47 0.0 201.61 0.07 ;
      LAYER M3 ;
      RECT 201.47 0.0 201.61 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[27]
  PIN TA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 383.16 0.0 383.3 0.07 ;
      LAYER M2 ;
      RECT 383.16 0.0 383.3 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[2]
  PIN TD[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 201.05 0.0 201.19 0.07 ;
      LAYER M3 ;
      RECT 201.05 0.0 201.19 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[27]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 383.41 0.0 383.55 0.07 ;
      LAYER M2 ;
      RECT 383.41 0.0 383.55 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[54]
  PIN DY[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 200.84 0.0 200.98 0.07 ;
      LAYER M1 ;
      RECT 200.84 0.0 200.98 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[27]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 383.98 0.0 384.12 0.07 ;
      LAYER M4 ;
      RECT 383.98 0.0 384.12 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[54]
  PIN TQ[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 199.5 0.0 199.64 0.07 ;
      LAYER M3 ;
      RECT 199.5 0.0 199.64 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[27]
  PIN TD[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 384.4 0.0 384.54 0.07 ;
      LAYER M4 ;
      RECT 384.4 0.0 384.54 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[54]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 195.4 0.0 195.54 0.07 ;
      LAYER M1 ;
      RECT 195.4 0.0 195.54 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[26]
  PIN DY[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 384.61 0.0 384.75 0.07 ;
      LAYER M2 ;
      RECT 384.61 0.0 384.75 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[54]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 194.83 0.0 194.97 0.07 ;
      LAYER M3 ;
      RECT 194.83 0.0 194.97 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[26]
  PIN TQ[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 385.95 0.0 386.09 0.07 ;
      LAYER M4 ;
      RECT 385.95 0.0 386.09 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[54]
  PIN TD[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 194.41 0.0 194.55 0.07 ;
      LAYER M3 ;
      RECT 194.41 0.0 194.55 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[26]
  PIN AY[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 386.215 0.0 386.355 0.07 ;
      LAYER M2 ;
      RECT 386.215 0.0 386.355 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[2]
  PIN DY[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 194.2 0.0 194.34 0.07 ;
      LAYER M1 ;
      RECT 194.2 0.0 194.34 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[26]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 387.195 0.0 387.335 0.07 ;
      LAYER M2 ;
      RECT 387.195 0.0 387.335 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[1]
  PIN TQ[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 192.86 0.0 193.0 0.07 ;
      LAYER M3 ;
      RECT 192.86 0.0 193.0 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[26]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 390.05 0.0 390.19 0.07 ;
      LAYER M2 ;
      RECT 390.05 0.0 390.19 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[55]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 188.76 0.0 188.9 0.07 ;
      LAYER M1 ;
      RECT 188.76 0.0 188.9 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[25]
  PIN TA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 390.3 0.0 390.44 0.07 ;
      LAYER M2 ;
      RECT 390.3 0.0 390.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[1]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 188.19 0.0 188.33 0.07 ;
      LAYER M3 ;
      RECT 188.19 0.0 188.33 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[25]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 390.62 0.0 390.76 0.07 ;
      LAYER M4 ;
      RECT 390.62 0.0 390.76 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[55]
  PIN TD[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 187.77 0.0 187.91 0.07 ;
      LAYER M3 ;
      RECT 187.77 0.0 187.91 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[25]
  PIN TD[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 391.04 0.0 391.18 0.07 ;
      LAYER M4 ;
      RECT 391.04 0.0 391.18 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[55]
  PIN DY[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 187.56 0.0 187.7 0.07 ;
      LAYER M1 ;
      RECT 187.56 0.0 187.7 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[25]
  PIN DY[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 391.25 0.0 391.39 0.07 ;
      LAYER M2 ;
      RECT 391.25 0.0 391.39 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[55]
  PIN TQ[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 186.22 0.0 186.36 0.07 ;
      LAYER M3 ;
      RECT 186.22 0.0 186.36 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[25]
  PIN TQ[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 392.59 0.0 392.73 0.07 ;
      LAYER M4 ;
      RECT 392.59 0.0 392.73 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[55]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 181.89 0.0 182.03 0.07 ;
      LAYER M1 ;
      RECT 181.89 0.0 182.03 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[24]
  PIN AY[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 392.945 0.0 393.085 0.07 ;
      LAYER M2 ;
      RECT 392.945 0.0 393.085 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[1]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 181.55 0.0 181.69 0.07 ;
      LAYER M3 ;
      RECT 181.55 0.0 181.69 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[24]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 393.785 0.0 393.925 0.07 ;
      LAYER M2 ;
      RECT 393.785 0.0 393.925 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END A[0]
  PIN TD[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 181.13 0.0 181.27 0.07 ;
      LAYER M3 ;
      RECT 181.13 0.0 181.27 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[24]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 396.69 0.0 396.83 0.07 ;
      LAYER M2 ;
      RECT 396.69 0.0 396.83 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[56]
  PIN DY[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 180.92 0.0 181.06 0.07 ;
      LAYER M1 ;
      RECT 180.92 0.0 181.06 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[24]
  PIN TA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 397.07 0.0 397.21 0.07 ;
      LAYER M2 ;
      RECT 397.07 0.0 397.21 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TA[0]
  PIN TQ[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 179.58 0.0 179.72 0.07 ;
      LAYER M3 ;
      RECT 179.58 0.0 179.72 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[24]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 397.26 0.0 397.4 0.07 ;
      LAYER M4 ;
      RECT 397.26 0.0 397.4 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[56]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 175.48 0.0 175.62 0.07 ;
      LAYER M1 ;
      RECT 175.48 0.0 175.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[23]
  PIN TD[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 397.68 0.0 397.82 0.07 ;
      LAYER M4 ;
      RECT 397.68 0.0 397.82 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[56]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 174.91 0.0 175.05 0.07 ;
      LAYER M3 ;
      RECT 174.91 0.0 175.05 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[23]
  PIN DY[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 397.89 0.0 398.03 0.07 ;
      LAYER M2 ;
      RECT 397.89 0.0 398.03 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[56]
  PIN TD[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 174.49 0.0 174.63 0.07 ;
      LAYER M3 ;
      RECT 174.49 0.0 174.63 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[23]
  PIN TQ[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 399.23 0.0 399.37 0.07 ;
      LAYER M4 ;
      RECT 399.23 0.0 399.37 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[56]
  PIN DY[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 174.28 0.0 174.42 0.07 ;
      LAYER M1 ;
      RECT 174.28 0.0 174.42 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[23]
  PIN AY[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 400.26 0.0 400.4 0.07 ;
      LAYER M2 ;
      RECT 400.26 0.0 400.4 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END AY[0]
  PIN TQ[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 172.94 0.0 173.08 0.07 ;
      LAYER M3 ;
      RECT 172.94 0.0 173.08 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[23]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 403.33 0.0 403.47 0.07 ;
      LAYER M2 ;
      RECT 403.33 0.0 403.47 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[57]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 168.84 0.0 168.98 0.07 ;
      LAYER M1 ;
      RECT 168.84 0.0 168.98 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[22]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 403.9 0.0 404.04 0.07 ;
      LAYER M4 ;
      RECT 403.9 0.0 404.04 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[57]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 168.27 0.0 168.41 0.07 ;
      LAYER M3 ;
      RECT 168.27 0.0 168.41 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[22]
  PIN TD[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 404.32 0.0 404.46 0.07 ;
      LAYER M4 ;
      RECT 404.32 0.0 404.46 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[57]
  PIN TD[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 167.85 0.0 167.99 0.07 ;
      LAYER M3 ;
      RECT 167.85 0.0 167.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[22]
  PIN DY[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 404.53 0.0 404.67 0.07 ;
      LAYER M2 ;
      RECT 404.53 0.0 404.67 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[57]
  PIN DY[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 167.64 0.0 167.78 0.07 ;
      LAYER M1 ;
      RECT 167.64 0.0 167.78 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[22]
  PIN TQ[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 405.87 0.0 406.01 0.07 ;
      LAYER M4 ;
      RECT 405.87 0.0 406.01 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[57]
  PIN TQ[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 166.3 0.0 166.44 0.07 ;
      LAYER M3 ;
      RECT 166.3 0.0 166.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[22]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 409.97 0.0 410.11 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[58]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 162.2 0.0 162.34 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[21]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 410.54 0.0 410.68 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[58]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 161.63 0.0 161.77 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[21]
  PIN TD[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 410.96 0.0 411.1 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[58]
  PIN TD[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 161.21 0.0 161.35 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[21]
  PIN DY[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 411.17 0.0 411.31 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[58]
  PIN DY[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 161.0 0.0 161.14 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[21]
  PIN TQ[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 412.51 0.0 412.65 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[58]
  PIN TQ[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 159.66 0.0 159.8 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[21]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 416.61 0.0 416.75 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[59]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 155.56 0.0 155.7 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[20]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 417.18 0.0 417.32 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[59]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 154.99 0.0 155.13 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[20]
  PIN TD[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 417.6 0.0 417.74 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[59]
  PIN TD[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 154.57 0.0 154.71 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[20]
  PIN DY[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 417.81 0.0 417.95 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[59]
  PIN DY[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 154.36 0.0 154.5 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[20]
  PIN TQ[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 419.15 0.0 419.29 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[59]
  PIN TQ[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 153.02 0.0 153.16 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[20]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 441.81 0.0 441.95 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[60]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 130.36 0.0 130.5 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[19]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 442.38 0.0 442.52 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[60]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 129.79 0.0 129.93 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[19]
  PIN TD[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 442.8 0.0 442.94 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[60]
  PIN TD[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 129.37 0.0 129.51 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[19]
  PIN DY[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 443.01 0.0 443.15 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[60]
  PIN DY[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 129.16 0.0 129.3 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[19]
  PIN TQ[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 444.35 0.0 444.49 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[60]
  PIN TQ[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 127.82 0.0 127.96 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[19]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 448.45 0.0 448.59 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[61]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 123.72 0.0 123.86 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[18]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 449.02 0.0 449.16 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[61]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 123.15 0.0 123.29 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[18]
  PIN TD[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 449.44 0.0 449.58 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[61]
  PIN TD[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 122.73 0.0 122.87 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[18]
  PIN DY[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 449.65 0.0 449.79 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[61]
  PIN DY[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 122.52 0.0 122.66 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[18]
  PIN TQ[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 450.99 0.0 451.13 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[61]
  PIN TQ[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 121.18 0.0 121.32 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[18]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 455.09 0.0 455.23 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[62]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 117.08 0.0 117.22 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[17]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 455.66 0.0 455.8 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[62]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 116.51 0.0 116.65 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[17]
  PIN TD[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 456.08 0.0 456.22 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[62]
  PIN TD[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 116.09 0.0 116.23 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[17]
  PIN DY[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 456.29 0.0 456.43 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[62]
  PIN DY[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 115.88 0.0 116.02 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[17]
  PIN TQ[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 457.63 0.0 457.77 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[62]
  PIN TQ[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 114.54 0.0 114.68 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[17]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 461.73 0.0 461.87 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[63]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 110.44 0.0 110.58 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[16]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 462.3 0.0 462.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[63]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 109.87 0.0 110.01 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[16]
  PIN TD[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 462.72 0.0 462.86 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[63]
  PIN TD[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 109.45 0.0 109.59 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[16]
  PIN DY[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 462.93 0.0 463.07 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[63]
  PIN DY[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 109.24 0.0 109.38 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[16]
  PIN TQ[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 464.27 0.0 464.41 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[63]
  PIN TQ[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 107.9 0.0 108.04 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[16]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 468.37 0.0 468.51 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[64]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 103.8 0.0 103.94 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[15]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 468.94 0.0 469.08 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[64]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 103.23 0.0 103.37 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[15]
  PIN TD[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 469.36 0.0 469.5 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[64]
  PIN TD[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 102.81 0.0 102.95 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[15]
  PIN DY[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 469.57 0.0 469.71 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[64]
  PIN DY[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 102.6 0.0 102.74 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[15]
  PIN TQ[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 470.91 0.0 471.05 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[64]
  PIN TQ[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 101.26 0.0 101.4 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[15]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 475.01 0.0 475.15 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[65]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 97.16 0.0 97.3 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[14]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 475.58 0.0 475.72 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[65]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 96.59 0.0 96.73 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[14]
  PIN TD[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 476.0 0.0 476.14 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[65]
  PIN TD[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 96.17 0.0 96.31 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[14]
  PIN DY[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 476.21 0.0 476.35 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[65]
  PIN DY[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 95.96 0.0 96.1 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[14]
  PIN TQ[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 477.55 0.0 477.69 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[65]
  PIN TQ[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 94.62 0.0 94.76 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[14]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 481.65 0.0 481.79 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[66]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 90.52 0.0 90.66 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[13]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 482.22 0.0 482.36 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[66]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 89.95 0.0 90.09 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[13]
  PIN TD[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 482.64 0.0 482.78 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[66]
  PIN TD[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 89.53 0.0 89.67 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[13]
  PIN DY[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 482.85 0.0 482.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[66]
  PIN DY[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 89.32 0.0 89.46 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[13]
  PIN TQ[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 484.19 0.0 484.33 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[66]
  PIN TQ[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 87.98 0.0 88.12 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[13]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 488.29 0.0 488.43 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[67]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 83.88 0.0 84.02 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[12]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 488.86 0.0 489.0 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[67]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 83.31 0.0 83.45 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[12]
  PIN TD[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 489.28 0.0 489.42 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[67]
  PIN TD[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 82.89 0.0 83.03 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[12]
  PIN DY[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 489.49 0.0 489.63 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[67]
  PIN DY[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 82.68 0.0 82.82 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[12]
  PIN TQ[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 490.83 0.0 490.97 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[67]
  PIN TQ[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 81.34 0.0 81.48 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[12]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 494.93 0.0 495.07 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[68]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 77.24 0.0 77.38 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[11]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 495.5 0.0 495.64 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[68]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 76.67 0.0 76.81 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[11]
  PIN TD[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 495.92 0.0 496.06 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[68]
  PIN TD[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 76.25 0.0 76.39 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[11]
  PIN DY[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 496.13 0.0 496.27 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[68]
  PIN DY[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 76.04 0.0 76.18 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[11]
  PIN TQ[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 497.47 0.0 497.61 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[68]
  PIN TQ[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 74.7 0.0 74.84 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[11]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 501.57 0.0 501.71 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[69]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 70.6 0.0 70.74 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[10]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 502.14 0.0 502.28 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[69]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 70.03 0.0 70.17 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[10]
  PIN TD[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 502.56 0.0 502.7 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[69]
  PIN TD[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 69.61 0.0 69.75 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[10]
  PIN DY[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 502.77 0.0 502.91 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[69]
  PIN DY[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 69.4 0.0 69.54 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[10]
  PIN TQ[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 504.11 0.0 504.25 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[69]
  PIN TQ[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 68.06 0.0 68.2 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[10]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 508.21 0.0 508.35 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[70]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 63.96 0.0 64.1 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[9]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 508.78 0.0 508.92 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[70]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 63.39 0.0 63.53 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[9]
  PIN TD[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 509.2 0.0 509.34 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[70]
  PIN TD[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 62.97 0.0 63.11 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[9]
  PIN DY[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 509.41 0.0 509.55 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[70]
  PIN DY[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 62.76 0.0 62.9 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[9]
  PIN TQ[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 510.75 0.0 510.89 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[70]
  PIN TQ[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 61.42 0.0 61.56 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[9]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 514.85 0.0 514.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[71]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 57.32 0.0 57.46 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[8]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 515.42 0.0 515.56 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[71]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 56.75 0.0 56.89 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[8]
  PIN TD[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 515.84 0.0 515.98 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[71]
  PIN TD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 56.33 0.0 56.47 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[8]
  PIN DY[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 516.05 0.0 516.19 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[71]
  PIN DY[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 56.12 0.0 56.26 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[8]
  PIN TQ[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 517.39 0.0 517.53 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[71]
  PIN TQ[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 54.78 0.0 54.92 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[8]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 521.49 0.0 521.63 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[72]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 50.68 0.0 50.82 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[7]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 522.06 0.0 522.2 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[72]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 50.11 0.0 50.25 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[7]
  PIN TD[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 522.48 0.0 522.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[72]
  PIN TD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 49.69 0.0 49.83 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[7]
  PIN DY[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 522.69 0.0 522.83 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[72]
  PIN DY[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 49.48 0.0 49.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[7]
  PIN TQ[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 524.03 0.0 524.17 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[72]
  PIN TQ[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 48.14 0.0 48.28 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[7]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 528.13 0.0 528.27 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[73]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 44.04 0.0 44.18 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[6]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 528.7 0.0 528.84 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[73]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 43.47 0.0 43.61 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[6]
  PIN TD[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 529.12 0.0 529.26 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[73]
  PIN TD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 43.05 0.0 43.19 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[6]
  PIN DY[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 529.33 0.0 529.47 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[73]
  PIN DY[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 42.84 0.0 42.98 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[6]
  PIN TQ[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 530.67 0.0 530.81 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[73]
  PIN TQ[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 41.5 0.0 41.64 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[6]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 534.77 0.0 534.91 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[74]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 37.4 0.0 37.54 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[5]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 535.34 0.0 535.48 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[74]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 36.83 0.0 36.97 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[5]
  PIN TD[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 535.76 0.0 535.9 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[74]
  PIN TD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 36.41 0.0 36.55 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[5]
  PIN DY[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 535.97 0.0 536.11 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[74]
  PIN DY[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 36.2 0.0 36.34 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[5]
  PIN TQ[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 537.31 0.0 537.45 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[74]
  PIN TQ[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 34.86 0.0 35.0 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[5]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 541.41 0.0 541.55 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[75]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 30.76 0.0 30.9 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[4]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 541.98 0.0 542.12 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[75]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 30.19 0.0 30.33 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[4]
  PIN TD[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 542.4 0.0 542.54 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[75]
  PIN TD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 29.77 0.0 29.91 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[4]
  PIN DY[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 542.61 0.0 542.75 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[75]
  PIN DY[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 29.56 0.0 29.7 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[4]
  PIN TQ[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 543.95 0.0 544.09 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[75]
  PIN TQ[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 28.22 0.0 28.36 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[4]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 548.05 0.0 548.19 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[76]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 24.12 0.0 24.26 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[3]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 548.62 0.0 548.76 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[76]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 23.55 0.0 23.69 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[3]
  PIN TD[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 549.04 0.0 549.18 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[76]
  PIN TD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 23.13 0.0 23.27 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[3]
  PIN DY[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 549.25 0.0 549.39 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[76]
  PIN DY[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 22.92 0.0 23.06 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[3]
  PIN TQ[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 550.59 0.0 550.73 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[76]
  PIN TQ[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 21.58 0.0 21.72 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[3]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 554.69 0.0 554.83 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[77]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 17.48 0.0 17.62 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[2]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 555.26 0.0 555.4 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[77]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.91 0.0 17.05 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[2]
  PIN TD[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 555.68 0.0 555.82 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[77]
  PIN TD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.49 0.0 16.63 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[2]
  PIN DY[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 555.89 0.0 556.03 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[77]
  PIN DY[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 16.28 0.0 16.42 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[2]
  PIN TQ[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 557.23 0.0 557.37 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[77]
  PIN TQ[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 14.94 0.0 15.08 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[2]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 561.33 0.0 561.47 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[78]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 10.84 0.0 10.98 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[1]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 561.9 0.0 562.04 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[78]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.27 0.0 10.41 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[1]
  PIN TD[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 562.32 0.0 562.46 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[78]
  PIN TD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 9.85 0.0 9.99 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[1]
  PIN DY[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 562.53 0.0 562.67 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[78]
  PIN DY[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 9.64 0.0 9.78 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[1]
  PIN TQ[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 563.87 0.0 564.01 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[78]
  PIN TQ[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 8.3 0.0 8.44 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[1]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 567.97 0.0 568.11 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[79]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 4.2 0.0 4.34 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END D[0]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 568.54 0.0 568.68 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[79]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 3.63 0.0 3.77 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END Q[0]
  PIN TD[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 568.96 0.0 569.1 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[79]
  PIN TD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 3.21 0.0 3.35 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TD[0]
  PIN DY[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 569.17 0.0 569.31 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[79]
  PIN DY[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 3.0 0.0 3.14 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END DY[0]
  PIN TQ[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 570.51 0.0 570.65 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[79]
  PIN TQ[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 1.66 0.0 1.8 0.07 ;
      END
    ANTENNAGATEAREA 0.0048 ;
    ANTENNADIFFAREA 0.06 ;
    END TQ[0]
  PIN VDDPE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 3.88 0.0 4.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.2 0.0 7.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.52 0.0 10.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 13.84 0.0 14.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.16 0.0 17.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.48 0.0 20.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 23.8 0.0 24.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.12 0.0 27.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.44 0.0 30.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 33.76 0.0 33.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.08 0.0 37.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 40.4 0.0 40.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 43.72 0.0 43.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.04 0.0 47.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.36 0.0 50.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 53.68 0.0 53.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 57.0 0.0 57.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 60.32 0.0 60.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 63.64 0.0 63.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 66.96 0.0 67.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.28 0.0 70.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 73.6 0.0 73.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 76.92 0.0 77.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 80.24 0.0 80.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 83.56 0.0 83.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 86.88 0.0 87.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.2 0.0 90.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 93.52 0.0 93.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 96.84 0.0 97.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.16 0.0 100.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.48 0.0 103.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 106.8 0.0 107.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 110.12 0.0 110.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 113.44 0.0 113.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 116.76 0.0 116.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.08 0.0 120.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.4 0.0 123.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 126.72 0.0 126.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 130.04 0.0 130.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 133.36 0.0 133.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.165 0.0 144.385 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 155.24 0.0 155.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 158.56 0.0 158.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 161.88 0.0 162.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 165.2 0.0 165.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 168.52 0.0 168.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 171.84 0.0 172.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 175.16 0.0 175.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 178.48 0.0 178.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 181.8 0.0 182.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 185.12 0.0 185.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 188.44 0.0 188.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 191.76 0.0 191.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 195.08 0.0 195.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 198.4 0.0 198.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 201.72 0.0 201.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 205.04 0.0 205.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 208.36 0.0 208.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 211.68 0.0 211.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.0 0.0 215.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 218.32 0.0 218.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 221.64 0.0 221.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 224.96 0.0 225.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 228.28 0.0 228.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 231.6 0.0 231.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 234.92 0.0 235.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 238.24 0.0 238.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 241.56 0.0 241.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 244.88 0.0 245.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 248.2 0.0 248.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 251.52 0.0 251.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 254.84 0.0 255.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 258.16 0.0 258.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 261.48 0.0 261.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 264.8 0.0 265.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 268.12 0.0 268.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 271.44 0.0 271.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 274.76 0.0 274.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 278.08 0.0 278.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 281.4 0.0 281.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 284.72 0.0 284.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 287.38 0.0 287.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 290.7 0.0 290.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 294.02 0.0 294.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 297.34 0.0 297.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 300.66 0.0 300.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 303.98 0.0 304.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 307.3 0.0 307.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 310.62 0.0 310.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 313.94 0.0 314.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 317.26 0.0 317.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 320.58 0.0 320.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 323.9 0.0 324.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 327.22 0.0 327.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 330.54 0.0 330.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 333.86 0.0 334.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 337.18 0.0 337.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 340.5 0.0 340.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 343.82 0.0 344.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 347.14 0.0 347.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 350.46 0.0 350.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 353.78 0.0 353.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 357.1 0.0 357.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 360.42 0.0 360.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 363.74 0.0 363.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 367.06 0.0 367.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 370.38 0.0 370.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 373.7 0.0 373.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 377.02 0.0 377.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 380.34 0.0 380.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 383.66 0.0 383.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 386.98 0.0 387.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 390.3 0.0 390.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 393.62 0.0 393.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 396.94 0.0 397.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 400.26 0.0 400.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 403.58 0.0 403.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 406.9 0.0 407.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 410.22 0.0 410.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 413.54 0.0 413.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 416.86 0.0 417.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 427.925 0.0 428.145 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 438.74 0.0 438.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 442.06 0.0 442.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 445.38 0.0 445.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 448.7 0.0 448.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 452.02 0.0 452.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 455.34 0.0 455.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 458.66 0.0 458.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 461.98 0.0 462.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 465.3 0.0 465.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 468.62 0.0 468.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 471.94 0.0 472.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 475.26 0.0 475.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 478.58 0.0 478.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 481.9 0.0 482.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 485.22 0.0 485.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 488.54 0.0 488.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 491.86 0.0 492.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 495.18 0.0 495.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 498.5 0.0 498.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 501.82 0.0 502.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 505.14 0.0 505.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 508.46 0.0 508.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 511.78 0.0 511.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 515.1 0.0 515.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 518.42 0.0 518.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 521.74 0.0 521.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 525.06 0.0 525.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 528.38 0.0 528.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 531.7 0.0 531.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 535.02 0.0 535.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 538.34 0.0 538.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 541.66 0.0 541.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 544.98 0.0 545.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 548.3 0.0 548.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 551.62 0.0 551.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 554.94 0.0 555.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 558.26 0.0 558.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 561.58 0.0 561.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 564.9 0.0 565.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 568.22 0.0 568.43 145.84 ;
      END
    END VDDPE
  PIN VDDCE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 1.34 0.0 1.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 4.66 0.0 4.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.98 0.0 8.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 11.3 0.0 11.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 14.62 0.0 14.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.94 0.0 18.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 21.26 0.0 21.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 24.58 0.0 24.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.9 0.0 28.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 31.22 0.0 31.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 34.54 0.0 34.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.86 0.0 38.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 41.18 0.0 41.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.5 0.0 44.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.82 0.0 48.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.14 0.0 51.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 54.46 0.0 54.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 57.78 0.0 57.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.1 0.0 61.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.42 0.0 64.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.74 0.0 67.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 71.06 0.0 71.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.38 0.0 74.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 77.7 0.0 77.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.02 0.0 81.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.34 0.0 84.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.66 0.0 87.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.98 0.0 91.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.3 0.0 94.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 97.62 0.0 97.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.94 0.0 101.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 104.26 0.0 104.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 107.58 0.0 107.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 110.9 0.0 111.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 114.22 0.0 114.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 117.54 0.0 117.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.86 0.0 121.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 124.18 0.0 124.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 127.5 0.0 127.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 130.82 0.0 131.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.595 0.0 147.815 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 152.7 0.0 152.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.02 0.0 156.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 159.34 0.0 159.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 162.66 0.0 162.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 165.98 0.0 166.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 169.3 0.0 169.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 172.62 0.0 172.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 175.94 0.0 176.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 179.26 0.0 179.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 182.58 0.0 182.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 185.9 0.0 186.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 189.22 0.0 189.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 192.54 0.0 192.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 195.86 0.0 196.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.18 0.0 199.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 202.5 0.0 202.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 205.82 0.0 206.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 209.14 0.0 209.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 212.46 0.0 212.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.78 0.0 215.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 219.1 0.0 219.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 222.42 0.0 222.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.74 0.0 225.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.06 0.0 229.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.38 0.0 232.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.7 0.0 235.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.02 0.0 239.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.34 0.0 242.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 245.66 0.0 245.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 248.98 0.0 249.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.3 0.0 252.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 255.62 0.0 255.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 258.94 0.0 259.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.26 0.0 262.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 265.58 0.0 265.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 268.9 0.0 269.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 272.22 0.0 272.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 275.54 0.0 275.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 278.86 0.0 279.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 282.18 0.0 282.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 289.92 0.0 290.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 293.24 0.0 293.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 296.56 0.0 296.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 299.88 0.0 300.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 303.2 0.0 303.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 306.52 0.0 306.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 309.84 0.0 310.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 313.16 0.0 313.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 316.48 0.0 316.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 319.8 0.0 320.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 323.12 0.0 323.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 326.44 0.0 326.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 329.76 0.0 329.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 333.08 0.0 333.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 336.4 0.0 336.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 339.72 0.0 339.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 343.04 0.0 343.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 346.36 0.0 346.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 349.68 0.0 349.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 353.0 0.0 353.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 356.32 0.0 356.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 359.64 0.0 359.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 362.96 0.0 363.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 366.28 0.0 366.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 369.6 0.0 369.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 372.92 0.0 373.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 376.24 0.0 376.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 379.56 0.0 379.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 382.88 0.0 383.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 386.2 0.0 386.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 389.52 0.0 389.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 392.84 0.0 393.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 396.16 0.0 396.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 399.48 0.0 399.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 402.8 0.0 403.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 406.12 0.0 406.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 409.44 0.0 409.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 412.76 0.0 412.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 416.08 0.0 416.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 419.4 0.0 419.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 424.495 0.0 424.715 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 441.28 0.0 441.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 444.6 0.0 444.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 447.92 0.0 448.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 451.24 0.0 451.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 454.56 0.0 454.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 457.88 0.0 458.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 461.2 0.0 461.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 464.52 0.0 464.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 467.84 0.0 468.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 471.16 0.0 471.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 474.48 0.0 474.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 477.8 0.0 478.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 481.12 0.0 481.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 484.44 0.0 484.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 487.76 0.0 487.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 491.08 0.0 491.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 494.4 0.0 494.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 497.72 0.0 497.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 501.04 0.0 501.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 504.36 0.0 504.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 507.68 0.0 507.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 511.0 0.0 511.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 514.32 0.0 514.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 517.64 0.0 517.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 520.96 0.0 521.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 524.28 0.0 524.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 527.6 0.0 527.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 530.92 0.0 531.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 534.24 0.0 534.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 537.56 0.0 537.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 540.88 0.0 541.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 544.2 0.0 544.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 547.52 0.0 547.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 550.84 0.0 551.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 554.16 0.0 554.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 557.48 0.0 557.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 560.8 0.0 561.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 564.12 0.0 564.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 567.44 0.0 567.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 570.76 0.0 570.97 145.84 ;
      END
    END VDDCE
  PIN VSSE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 2.68 0.0 2.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 6.0 0.0 6.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 9.32 0.0 9.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.64 0.0 12.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.96 0.0 16.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.28 0.0 19.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 22.6 0.0 22.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.92 0.0 26.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 29.24 0.0 29.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.56 0.0 32.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.88 0.0 36.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 39.2 0.0 39.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.52 0.0 42.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.84 0.0 46.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 49.16 0.0 49.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 52.48 0.0 52.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.8 0.0 56.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 59.12 0.0 59.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 62.44 0.0 62.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 65.76 0.0 65.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 69.08 0.0 69.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.4 0.0 72.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.72 0.0 75.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 79.04 0.0 79.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.36 0.0 82.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 85.68 0.0 85.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 89.0 0.0 89.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.32 0.0 92.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 95.64 0.0 95.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.96 0.0 99.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 102.28 0.0 102.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 105.6 0.0 105.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.92 0.0 109.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 112.24 0.0 112.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 115.56 0.0 115.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.88 0.0 119.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 122.2 0.0 122.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 125.52 0.0 125.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.84 0.0 129.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 132.16 0.0 132.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.845 0.0 145.065 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 154.04 0.0 154.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 157.36 0.0 157.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 160.68 0.0 160.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 164.0 0.0 164.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 167.32 0.0 167.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 170.64 0.0 170.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 173.96 0.0 174.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.28 0.0 177.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 180.6 0.0 180.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 183.92 0.0 184.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.24 0.0 187.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.56 0.0 190.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 193.88 0.0 194.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 197.2 0.0 197.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 200.52 0.0 200.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 203.84 0.0 204.05 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.16 0.0 207.37 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 210.48 0.0 210.69 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.8 0.0 214.01 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 217.12 0.0 217.33 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 220.44 0.0 220.65 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 223.76 0.0 223.97 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 227.08 0.0 227.29 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 230.4 0.0 230.61 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 233.72 0.0 233.93 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 237.04 0.0 237.25 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 240.36 0.0 240.57 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 243.68 0.0 243.89 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 247.0 0.0 247.21 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 250.32 0.0 250.53 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 253.64 0.0 253.85 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 256.96 0.0 257.17 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 260.28 0.0 260.49 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 263.6 0.0 263.81 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 266.92 0.0 267.13 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 270.24 0.0 270.45 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 273.56 0.0 273.77 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 276.88 0.0 277.09 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 280.2 0.0 280.41 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 283.52 0.0 283.73 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 288.58 0.0 288.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 291.9 0.0 292.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 295.22 0.0 295.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 298.54 0.0 298.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 301.86 0.0 302.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 305.18 0.0 305.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 308.5 0.0 308.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 311.82 0.0 312.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 315.14 0.0 315.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 318.46 0.0 318.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 321.78 0.0 321.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 325.1 0.0 325.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 328.42 0.0 328.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 331.74 0.0 331.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 335.06 0.0 335.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 338.38 0.0 338.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 341.7 0.0 341.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 345.02 0.0 345.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 348.34 0.0 348.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 351.66 0.0 351.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 354.98 0.0 355.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 358.3 0.0 358.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 361.62 0.0 361.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 364.94 0.0 365.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 368.26 0.0 368.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 371.58 0.0 371.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 374.9 0.0 375.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 378.22 0.0 378.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 381.54 0.0 381.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 384.86 0.0 385.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 388.18 0.0 388.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 391.5 0.0 391.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 394.82 0.0 395.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 398.14 0.0 398.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 401.46 0.0 401.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 404.78 0.0 404.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 408.1 0.0 408.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 411.42 0.0 411.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 414.74 0.0 414.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 418.06 0.0 418.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 427.245 0.0 427.465 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 439.94 0.0 440.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 443.26 0.0 443.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 446.58 0.0 446.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 449.9 0.0 450.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 453.22 0.0 453.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 456.54 0.0 456.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 459.86 0.0 460.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 463.18 0.0 463.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 466.5 0.0 466.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 469.82 0.0 470.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 473.14 0.0 473.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 476.46 0.0 476.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 479.78 0.0 479.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 483.1 0.0 483.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 486.42 0.0 486.63 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 489.74 0.0 489.95 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 493.06 0.0 493.27 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 496.38 0.0 496.59 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 499.7 0.0 499.91 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 503.02 0.0 503.23 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 506.34 0.0 506.55 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 509.66 0.0 509.87 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 512.98 0.0 513.19 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 516.3 0.0 516.51 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 519.62 0.0 519.83 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 522.94 0.0 523.15 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 526.26 0.0 526.47 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 529.58 0.0 529.79 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 532.9 0.0 533.11 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 536.22 0.0 536.43 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 539.54 0.0 539.75 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 542.86 0.0 543.07 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 546.18 0.0 546.39 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 549.5 0.0 549.71 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 552.82 0.0 553.03 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 556.14 0.0 556.35 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 559.46 0.0 559.67 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 562.78 0.0 562.99 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 566.1 0.0 566.31 145.84 ;
      END
    PORT
      LAYER M4 ;
      RECT 569.42 0.0 569.63 145.84 ;
      END
    END VSSE
  OBS
    #otc obstructions
    LAYER M1 DESIGNRULEWIDTH 0.07 ;
    RECT 404.74 0.0 572.31 0.14 ;
    RECT 403.54 0.0 404.46 0.14 ;
    RECT 400.47 0.0 403.26 0.14 ;
    RECT 398.1 0.0 400.19 0.14 ;
    RECT 397.28 0.0 397.82 0.14 ;
    RECT 396.9 0.0 397.0 0.14 ;
    RECT 393.995 0.0 396.62 0.14 ;
    RECT 393.155 0.0 393.715 0.14 ;
    RECT 391.46 0.0 392.875 0.14 ;
    RECT 390.51 0.0 391.18 0.14 ;
    RECT 387.405 0.0 389.98 0.14 ;
    RECT 386.425 0.0 387.125 0.14 ;
    RECT 384.82 0.0 386.145 0.14 ;
    RECT 383.62 0.0 384.54 0.14 ;
    RECT 379.74 0.0 383.09 0.14 ;
    RECT 378.18 0.0 379.46 0.14 ;
    RECT 376.98 0.0 377.9 0.14 ;
    RECT 371.54 0.0 376.7 0.14 ;
    RECT 370.34 0.0 371.26 0.14 ;
    RECT 364.9 0.0 370.06 0.14 ;
    RECT 364.115 0.0 364.62 0.14 ;
    RECT 363.7 0.0 363.835 0.14 ;
    RECT 362.605 0.0 363.42 0.14 ;
    RECT 359.285 0.0 362.325 0.14 ;
    RECT 358.58 0.0 359.005 0.14 ;
    RECT 357.06 0.0 357.98 0.14 ;
    RECT 353.165 0.0 356.78 0.14 ;
    RECT 352.645 0.0 352.885 0.14 ;
    RECT 351.975 0.0 352.365 0.14 ;
    RECT 350.42 0.0 351.34 0.14 ;
    RECT 346.005 0.0 350.14 0.14 ;
    RECT 345.335 0.0 345.725 0.14 ;
    RECT 343.78 0.0 344.7 0.14 ;
    RECT 338.34 0.0 343.5 0.14 ;
    RECT 337.14 0.0 338.06 0.14 ;
    RECT 331.7 0.0 336.86 0.14 ;
    RECT 330.5 0.0 331.42 0.14 ;
    RECT 327.535 0.0 330.22 0.14 ;
    RECT 325.06 0.0 327.255 0.14 ;
    RECT 324.39 0.0 324.78 0.14 ;
    RECT 323.86 0.0 324.11 0.14 ;
    RECT 322.06 0.0 323.58 0.14 ;
    RECT 320.29 0.0 321.78 0.14 ;
    RECT 319.45 0.0 320.01 0.14 ;
    RECT 318.42 0.0 319.17 0.14 ;
    RECT 317.22 0.0 318.14 0.14 ;
    RECT 314.315 0.0 316.94 0.14 ;
    RECT 313.405 0.0 314.035 0.14 ;
    RECT 311.78 0.0 313.125 0.14 ;
    RECT 310.995 0.0 311.5 0.14 ;
    RECT 310.58 0.0 310.715 0.14 ;
    RECT 307.51 0.0 310.3 0.14 ;
    RECT 306.745 0.0 307.23 0.14 ;
    RECT 305.14 0.0 306.465 0.14 ;
    RECT 303.94 0.0 304.86 0.14 ;
    RECT 301.035 0.0 303.41 0.14 ;
    RECT 298.82 0.0 300.755 0.14 ;
    RECT 297.55 0.0 298.22 0.14 ;
    RECT 294.415 0.0 297.02 0.14 ;
    RECT 292.215 0.0 294.135 0.14 ;
    RECT 291.02 0.0 291.58 0.14 ;
    RECT 286.505 0.0 290.38 0.14 ;
    RECT 283.48 0.0 285.615 0.14 ;
    RECT 282.425 0.0 283.2 0.14 ;
    RECT 281.19 0.0 282.145 0.14 ;
    RECT 279.14 0.0 280.91 0.14 ;
    RECT 278.445 0.0 278.86 0.14 ;
    RECT 275.655 0.0 278.165 0.14 ;
    RECT 274.51 0.0 275.375 0.14 ;
    RECT 269.015 0.0 274.23 0.14 ;
    RECT 267.87 0.0 268.735 0.14 ;
    RECT 266.35 0.0 267.59 0.14 ;
    RECT 264.09 0.0 266.07 0.14 ;
    RECT 262.375 0.0 263.81 0.14 ;
    RECT 261.23 0.0 262.095 0.14 ;
    RECT 259.75 0.0 260.95 0.14 ;
    RECT 255.735 0.0 259.47 0.14 ;
    RECT 254.17 0.0 255.455 0.14 ;
    RECT 252.0 0.0 253.89 0.14 ;
    RECT 248.73 0.0 251.72 0.14 ;
    RECT 247.53 0.0 248.45 0.14 ;
    RECT 243.675 0.0 247.25 0.14 ;
    RECT 242.09 0.0 243.395 0.14 ;
    RECT 240.89 0.0 241.81 0.14 ;
    RECT 239.86 0.0 240.61 0.14 ;
    RECT 235.45 0.0 239.58 0.14 ;
    RECT 234.25 0.0 235.17 0.14 ;
    RECT 230.645 0.0 233.97 0.14 ;
    RECT 228.81 0.0 230.365 0.14 ;
    RECT 227.61 0.0 228.53 0.14 ;
    RECT 225.205 0.0 227.33 0.14 ;
    RECT 222.17 0.0 224.925 0.14 ;
    RECT 220.97 0.0 221.89 0.14 ;
    RECT 219.84 0.0 220.69 0.14 ;
    RECT 215.53 0.0 219.56 0.14 ;
    RECT 214.33 0.0 215.25 0.14 ;
    RECT 208.89 0.0 214.05 0.14 ;
    RECT 207.69 0.0 208.61 0.14 ;
    RECT 202.25 0.0 207.41 0.14 ;
    RECT 201.05 0.0 201.97 0.14 ;
    RECT 195.61 0.0 200.77 0.14 ;
    RECT 194.41 0.0 195.33 0.14 ;
    RECT 188.97 0.0 194.13 0.14 ;
    RECT 187.77 0.0 188.69 0.14 ;
    RECT 182.1 0.0 187.49 0.14 ;
    RECT 181.13 0.0 181.82 0.14 ;
    RECT 175.69 0.0 180.85 0.14 ;
    RECT 174.49 0.0 175.41 0.14 ;
    RECT 169.05 0.0 174.21 0.14 ;
    RECT 167.85 0.0 168.77 0.14 ;
    RECT 0.0 0.0 167.57 0.14 ;
    RECT 0.0 0.14 572.31 145.84 ;
    LAYER VIA1 ;
    RECT 0.0 0.0 572.31 145.84 ;
    LAYER M2 DESIGNRULEWIDTH 0.07 ;
    RECT 569.38 0.0 572.31 0.14 ;
    RECT 568.18 0.0 569.1 0.14 ;
    RECT 562.74 0.0 567.9 0.14 ;
    RECT 561.54 0.0 562.46 0.14 ;
    RECT 556.1 0.0 561.26 0.14 ;
    RECT 554.9 0.0 555.82 0.14 ;
    RECT 549.46 0.0 554.62 0.14 ;
    RECT 548.26 0.0 549.18 0.14 ;
    RECT 542.82 0.0 547.98 0.14 ;
    RECT 541.62 0.0 542.54 0.14 ;
    RECT 536.18 0.0 541.34 0.14 ;
    RECT 534.98 0.0 535.9 0.14 ;
    RECT 529.54 0.0 534.7 0.14 ;
    RECT 528.34 0.0 529.26 0.14 ;
    RECT 522.9 0.0 528.06 0.14 ;
    RECT 521.7 0.0 522.62 0.14 ;
    RECT 516.26 0.0 521.42 0.14 ;
    RECT 515.06 0.0 515.98 0.14 ;
    RECT 509.62 0.0 514.78 0.14 ;
    RECT 508.42 0.0 509.34 0.14 ;
    RECT 502.98 0.0 508.14 0.14 ;
    RECT 501.78 0.0 502.7 0.14 ;
    RECT 496.34 0.0 501.5 0.14 ;
    RECT 495.14 0.0 496.06 0.14 ;
    RECT 489.7 0.0 494.86 0.14 ;
    RECT 488.5 0.0 489.42 0.14 ;
    RECT 483.06 0.0 488.22 0.14 ;
    RECT 481.86 0.0 482.78 0.14 ;
    RECT 476.42 0.0 481.58 0.14 ;
    RECT 475.22 0.0 476.14 0.14 ;
    RECT 469.78 0.0 474.94 0.14 ;
    RECT 468.58 0.0 469.5 0.14 ;
    RECT 463.14 0.0 468.3 0.14 ;
    RECT 461.94 0.0 462.86 0.14 ;
    RECT 456.5 0.0 461.66 0.14 ;
    RECT 455.3 0.0 456.22 0.14 ;
    RECT 449.86 0.0 455.02 0.14 ;
    RECT 448.66 0.0 449.58 0.14 ;
    RECT 443.22 0.0 448.38 0.14 ;
    RECT 442.02 0.0 442.94 0.14 ;
    RECT 418.02 0.0 441.74 0.14 ;
    RECT 416.82 0.0 417.74 0.14 ;
    RECT 411.38 0.0 416.54 0.14 ;
    RECT 410.18 0.0 411.1 0.14 ;
    RECT 404.74 0.0 409.9 0.14 ;
    RECT 403.54 0.0 404.46 0.14 ;
    RECT 400.47 0.0 403.26 0.14 ;
    RECT 398.1 0.0 400.19 0.14 ;
    RECT 397.28 0.0 397.82 0.14 ;
    RECT 396.9 0.0 397.0 0.14 ;
    RECT 393.995 0.0 396.62 0.14 ;
    RECT 393.155 0.0 393.715 0.14 ;
    RECT 391.46 0.0 392.875 0.14 ;
    RECT 390.51 0.0 391.18 0.14 ;
    RECT 387.405 0.0 389.98 0.14 ;
    RECT 386.425 0.0 387.125 0.14 ;
    RECT 384.82 0.0 386.145 0.14 ;
    RECT 383.62 0.0 384.54 0.14 ;
    RECT 379.74 0.0 383.09 0.14 ;
    RECT 378.18 0.0 379.46 0.14 ;
    RECT 376.98 0.0 377.9 0.14 ;
    RECT 371.54 0.0 376.7 0.14 ;
    RECT 370.34 0.0 371.26 0.14 ;
    RECT 364.9 0.0 370.06 0.14 ;
    RECT 364.115 0.0 364.62 0.14 ;
    RECT 363.7 0.0 363.835 0.14 ;
    RECT 362.605 0.0 363.42 0.14 ;
    RECT 359.285 0.0 362.325 0.14 ;
    RECT 358.58 0.0 359.005 0.14 ;
    RECT 357.06 0.0 357.98 0.14 ;
    RECT 353.165 0.0 356.78 0.14 ;
    RECT 352.645 0.0 352.885 0.14 ;
    RECT 351.975 0.0 352.365 0.14 ;
    RECT 350.42 0.0 351.34 0.14 ;
    RECT 346.005 0.0 350.14 0.14 ;
    RECT 345.335 0.0 345.725 0.14 ;
    RECT 343.78 0.0 344.7 0.14 ;
    RECT 338.34 0.0 343.5 0.14 ;
    RECT 337.14 0.0 338.06 0.14 ;
    RECT 331.7 0.0 336.86 0.14 ;
    RECT 330.5 0.0 331.42 0.14 ;
    RECT 327.535 0.0 330.22 0.14 ;
    RECT 325.06 0.0 327.255 0.14 ;
    RECT 324.39 0.0 324.78 0.14 ;
    RECT 323.86 0.0 324.11 0.14 ;
    RECT 322.06 0.0 323.58 0.14 ;
    RECT 320.29 0.0 321.78 0.14 ;
    RECT 319.45 0.0 320.01 0.14 ;
    RECT 318.42 0.0 319.17 0.14 ;
    RECT 317.22 0.0 318.14 0.14 ;
    RECT 314.315 0.0 316.94 0.14 ;
    RECT 313.405 0.0 314.035 0.14 ;
    RECT 311.78 0.0 313.125 0.14 ;
    RECT 310.995 0.0 311.5 0.14 ;
    RECT 310.58 0.0 310.715 0.14 ;
    RECT 307.51 0.0 310.3 0.14 ;
    RECT 306.745 0.0 307.23 0.14 ;
    RECT 305.14 0.0 306.465 0.14 ;
    RECT 303.94 0.0 304.86 0.14 ;
    RECT 301.035 0.0 303.41 0.14 ;
    RECT 298.82 0.0 300.755 0.14 ;
    RECT 297.55 0.0 298.22 0.14 ;
    RECT 294.415 0.0 297.02 0.14 ;
    RECT 292.215 0.0 294.135 0.14 ;
    RECT 291.02 0.0 291.58 0.14 ;
    RECT 286.505 0.0 290.38 0.14 ;
    RECT 283.48 0.0 285.615 0.14 ;
    RECT 282.425 0.0 283.2 0.14 ;
    RECT 281.19 0.0 282.145 0.14 ;
    RECT 279.14 0.0 280.91 0.14 ;
    RECT 278.445 0.0 278.86 0.14 ;
    RECT 275.655 0.0 278.165 0.14 ;
    RECT 274.51 0.0 275.375 0.14 ;
    RECT 269.015 0.0 274.23 0.14 ;
    RECT 267.87 0.0 268.735 0.14 ;
    RECT 266.35 0.0 267.59 0.14 ;
    RECT 264.09 0.0 266.07 0.14 ;
    RECT 262.375 0.0 263.81 0.14 ;
    RECT 261.23 0.0 262.095 0.14 ;
    RECT 259.75 0.0 260.95 0.14 ;
    RECT 255.735 0.0 259.47 0.14 ;
    RECT 254.17 0.0 255.455 0.14 ;
    RECT 252.0 0.0 253.89 0.14 ;
    RECT 248.73 0.0 251.72 0.14 ;
    RECT 247.53 0.0 248.45 0.14 ;
    RECT 243.675 0.0 247.25 0.14 ;
    RECT 242.09 0.0 243.395 0.14 ;
    RECT 240.89 0.0 241.81 0.14 ;
    RECT 239.86 0.0 240.61 0.14 ;
    RECT 235.45 0.0 239.58 0.14 ;
    RECT 234.25 0.0 235.17 0.14 ;
    RECT 230.645 0.0 233.97 0.14 ;
    RECT 228.81 0.0 230.365 0.14 ;
    RECT 227.61 0.0 228.53 0.14 ;
    RECT 225.205 0.0 227.33 0.14 ;
    RECT 222.17 0.0 224.925 0.14 ;
    RECT 220.97 0.0 221.89 0.14 ;
    RECT 219.84 0.0 220.69 0.14 ;
    RECT 215.53 0.0 219.56 0.14 ;
    RECT 214.33 0.0 215.25 0.14 ;
    RECT 208.89 0.0 214.05 0.14 ;
    RECT 207.69 0.0 208.61 0.14 ;
    RECT 202.25 0.0 207.41 0.14 ;
    RECT 201.05 0.0 201.97 0.14 ;
    RECT 195.61 0.0 200.77 0.14 ;
    RECT 194.41 0.0 195.33 0.14 ;
    RECT 188.97 0.0 194.13 0.14 ;
    RECT 187.77 0.0 188.69 0.14 ;
    RECT 182.1 0.0 187.49 0.14 ;
    RECT 181.13 0.0 181.82 0.14 ;
    RECT 175.69 0.0 180.85 0.14 ;
    RECT 174.49 0.0 175.41 0.14 ;
    RECT 169.05 0.0 174.21 0.14 ;
    RECT 167.85 0.0 168.77 0.14 ;
    RECT 162.41 0.0 167.57 0.14 ;
    RECT 161.21 0.0 162.13 0.14 ;
    RECT 155.77 0.0 160.93 0.14 ;
    RECT 154.57 0.0 155.49 0.14 ;
    RECT 130.57 0.0 154.29 0.14 ;
    RECT 129.37 0.0 130.29 0.14 ;
    RECT 123.93 0.0 129.09 0.14 ;
    RECT 122.73 0.0 123.65 0.14 ;
    RECT 117.29 0.0 122.45 0.14 ;
    RECT 116.09 0.0 117.01 0.14 ;
    RECT 110.65 0.0 115.81 0.14 ;
    RECT 109.45 0.0 110.37 0.14 ;
    RECT 104.01 0.0 109.17 0.14 ;
    RECT 102.81 0.0 103.73 0.14 ;
    RECT 97.37 0.0 102.53 0.14 ;
    RECT 96.17 0.0 97.09 0.14 ;
    RECT 90.73 0.0 95.89 0.14 ;
    RECT 89.53 0.0 90.45 0.14 ;
    RECT 84.09 0.0 89.25 0.14 ;
    RECT 82.89 0.0 83.81 0.14 ;
    RECT 77.45 0.0 82.61 0.14 ;
    RECT 76.25 0.0 77.17 0.14 ;
    RECT 70.81 0.0 75.97 0.14 ;
    RECT 69.61 0.0 70.53 0.14 ;
    RECT 64.17 0.0 69.33 0.14 ;
    RECT 62.97 0.0 63.89 0.14 ;
    RECT 57.53 0.0 62.69 0.14 ;
    RECT 56.33 0.0 57.25 0.14 ;
    RECT 50.89 0.0 56.05 0.14 ;
    RECT 49.69 0.0 50.61 0.14 ;
    RECT 44.25 0.0 49.41 0.14 ;
    RECT 43.05 0.0 43.97 0.14 ;
    RECT 37.61 0.0 42.77 0.14 ;
    RECT 36.41 0.0 37.33 0.14 ;
    RECT 30.97 0.0 36.13 0.14 ;
    RECT 29.77 0.0 30.69 0.14 ;
    RECT 24.33 0.0 29.49 0.14 ;
    RECT 23.13 0.0 24.05 0.14 ;
    RECT 17.69 0.0 22.85 0.14 ;
    RECT 16.49 0.0 17.41 0.14 ;
    RECT 11.05 0.0 16.21 0.14 ;
    RECT 9.85 0.0 10.77 0.14 ;
    RECT 4.41 0.0 9.57 0.14 ;
    RECT 3.21 0.0 4.13 0.14 ;
    RECT 0.0 0.0 2.93 0.14 ;
    RECT 0.0 0.14 572.31 145.84 ;
    LAYER VIA2 ;
    RECT 0.0 0.0 572.31 145.84 ;
    LAYER M3 DESIGNRULEWIDTH 0.07 ;
    RECT 406.08 0.0 572.31 0.14 ;
    RECT 404.53 0.0 405.8 0.14 ;
    RECT 404.11 0.0 404.25 0.14 ;
    RECT 399.44 0.0 403.83 0.14 ;
    RECT 397.89 0.0 399.16 0.14 ;
    RECT 397.47 0.0 397.61 0.14 ;
    RECT 392.8 0.0 397.19 0.14 ;
    RECT 391.25 0.0 392.52 0.14 ;
    RECT 390.83 0.0 390.97 0.14 ;
    RECT 386.16 0.0 390.55 0.14 ;
    RECT 384.61 0.0 385.88 0.14 ;
    RECT 384.19 0.0 384.33 0.14 ;
    RECT 379.52 0.0 383.91 0.14 ;
    RECT 377.97 0.0 379.24 0.14 ;
    RECT 377.55 0.0 377.69 0.14 ;
    RECT 372.88 0.0 377.27 0.14 ;
    RECT 371.33 0.0 372.6 0.14 ;
    RECT 370.91 0.0 371.05 0.14 ;
    RECT 366.24 0.0 370.63 0.14 ;
    RECT 364.69 0.0 365.96 0.14 ;
    RECT 364.27 0.0 364.41 0.14 ;
    RECT 359.6 0.0 363.99 0.14 ;
    RECT 358.05 0.0 359.32 0.14 ;
    RECT 357.63 0.0 357.77 0.14 ;
    RECT 352.96 0.0 357.35 0.14 ;
    RECT 351.41 0.0 352.68 0.14 ;
    RECT 350.99 0.0 351.13 0.14 ;
    RECT 346.32 0.0 350.71 0.14 ;
    RECT 344.77 0.0 346.04 0.14 ;
    RECT 344.35 0.0 344.49 0.14 ;
    RECT 339.68 0.0 344.07 0.14 ;
    RECT 338.13 0.0 339.4 0.14 ;
    RECT 337.71 0.0 337.85 0.14 ;
    RECT 333.04 0.0 337.43 0.14 ;
    RECT 331.49 0.0 332.76 0.14 ;
    RECT 331.07 0.0 331.21 0.14 ;
    RECT 326.4 0.0 330.79 0.14 ;
    RECT 324.85 0.0 326.12 0.14 ;
    RECT 324.43 0.0 324.57 0.14 ;
    RECT 319.76 0.0 324.15 0.14 ;
    RECT 318.21 0.0 319.48 0.14 ;
    RECT 317.79 0.0 317.93 0.14 ;
    RECT 313.12 0.0 317.51 0.14 ;
    RECT 311.57 0.0 312.84 0.14 ;
    RECT 311.15 0.0 311.29 0.14 ;
    RECT 306.48 0.0 310.87 0.14 ;
    RECT 304.93 0.0 306.2 0.14 ;
    RECT 304.51 0.0 304.65 0.14 ;
    RECT 299.84 0.0 304.23 0.14 ;
    RECT 298.29 0.0 299.56 0.14 ;
    RECT 297.87 0.0 298.01 0.14 ;
    RECT 293.2 0.0 297.59 0.14 ;
    RECT 291.65 0.0 292.92 0.14 ;
    RECT 291.23 0.0 291.37 0.14 ;
    RECT 281.36 0.0 290.95 0.14 ;
    RECT 280.94 0.0 281.08 0.14 ;
    RECT 279.39 0.0 280.66 0.14 ;
    RECT 274.72 0.0 279.11 0.14 ;
    RECT 274.3 0.0 274.44 0.14 ;
    RECT 272.75 0.0 274.02 0.14 ;
    RECT 268.08 0.0 272.47 0.14 ;
    RECT 267.66 0.0 267.8 0.14 ;
    RECT 266.11 0.0 267.38 0.14 ;
    RECT 261.44 0.0 265.83 0.14 ;
    RECT 261.02 0.0 261.16 0.14 ;
    RECT 259.47 0.0 260.74 0.14 ;
    RECT 254.8 0.0 259.19 0.14 ;
    RECT 254.38 0.0 254.52 0.14 ;
    RECT 252.83 0.0 254.1 0.14 ;
    RECT 248.16 0.0 252.55 0.14 ;
    RECT 247.74 0.0 247.88 0.14 ;
    RECT 246.19 0.0 247.46 0.14 ;
    RECT 241.52 0.0 245.91 0.14 ;
    RECT 241.1 0.0 241.24 0.14 ;
    RECT 239.55 0.0 240.82 0.14 ;
    RECT 234.88 0.0 239.27 0.14 ;
    RECT 234.46 0.0 234.6 0.14 ;
    RECT 232.91 0.0 234.18 0.14 ;
    RECT 228.24 0.0 232.63 0.14 ;
    RECT 227.82 0.0 227.96 0.14 ;
    RECT 226.27 0.0 227.54 0.14 ;
    RECT 221.6 0.0 225.99 0.14 ;
    RECT 221.18 0.0 221.32 0.14 ;
    RECT 219.63 0.0 220.9 0.14 ;
    RECT 214.96 0.0 219.35 0.14 ;
    RECT 214.54 0.0 214.68 0.14 ;
    RECT 212.99 0.0 214.26 0.14 ;
    RECT 208.32 0.0 212.71 0.14 ;
    RECT 207.9 0.0 208.04 0.14 ;
    RECT 206.35 0.0 207.62 0.14 ;
    RECT 201.68 0.0 206.07 0.14 ;
    RECT 201.26 0.0 201.4 0.14 ;
    RECT 199.71 0.0 200.98 0.14 ;
    RECT 195.04 0.0 199.43 0.14 ;
    RECT 194.62 0.0 194.76 0.14 ;
    RECT 193.07 0.0 194.34 0.14 ;
    RECT 188.4 0.0 192.79 0.14 ;
    RECT 187.98 0.0 188.12 0.14 ;
    RECT 186.43 0.0 187.7 0.14 ;
    RECT 181.76 0.0 186.15 0.14 ;
    RECT 181.34 0.0 181.48 0.14 ;
    RECT 179.79 0.0 181.06 0.14 ;
    RECT 175.12 0.0 179.51 0.14 ;
    RECT 174.7 0.0 174.84 0.14 ;
    RECT 173.15 0.0 174.42 0.14 ;
    RECT 168.48 0.0 172.87 0.14 ;
    RECT 168.06 0.0 168.2 0.14 ;
    RECT 166.51 0.0 167.78 0.14 ;
    RECT 0.0 0.0 166.23 0.14 ;
    RECT 0.0 0.14 572.31 145.84 ;
    LAYER VIA3 ;
    RECT 0.0 0.0 572.31 145.84 ;
    LAYER M4 DESIGNRULEWIDTH 0.07 ;
    RECT 571.04 0.0 572.31 0.14 ;
    RECT 569.7 0.0 570.44 0.14 ;
    RECT 569.17 0.0 569.35 0.14 ;
    RECT 568.75 0.0 568.89 0.14 ;
    RECT 567.72 0.0 568.15 0.14 ;
    RECT 566.38 0.0 567.37 0.14 ;
    RECT 565.18 0.0 566.03 0.14 ;
    RECT 564.4 0.0 564.83 0.14 ;
    RECT 563.06 0.0 563.8 0.14 ;
    RECT 562.53 0.0 562.71 0.14 ;
    RECT 562.11 0.0 562.25 0.14 ;
    RECT 561.08 0.0 561.51 0.14 ;
    RECT 559.74 0.0 560.73 0.14 ;
    RECT 558.54 0.0 559.39 0.14 ;
    RECT 557.76 0.0 558.19 0.14 ;
    RECT 556.42 0.0 557.16 0.14 ;
    RECT 555.89 0.0 556.07 0.14 ;
    RECT 555.47 0.0 555.61 0.14 ;
    RECT 554.44 0.0 554.87 0.14 ;
    RECT 553.1 0.0 554.09 0.14 ;
    RECT 551.9 0.0 552.75 0.14 ;
    RECT 551.12 0.0 551.55 0.14 ;
    RECT 549.78 0.0 550.52 0.14 ;
    RECT 549.25 0.0 549.43 0.14 ;
    RECT 548.83 0.0 548.97 0.14 ;
    RECT 547.8 0.0 548.23 0.14 ;
    RECT 546.46 0.0 547.45 0.14 ;
    RECT 545.26 0.0 546.11 0.14 ;
    RECT 544.48 0.0 544.91 0.14 ;
    RECT 543.14 0.0 543.88 0.14 ;
    RECT 542.61 0.0 542.79 0.14 ;
    RECT 542.19 0.0 542.33 0.14 ;
    RECT 541.16 0.0 541.59 0.14 ;
    RECT 539.82 0.0 540.81 0.14 ;
    RECT 538.62 0.0 539.47 0.14 ;
    RECT 537.84 0.0 538.27 0.14 ;
    RECT 536.5 0.0 537.24 0.14 ;
    RECT 535.97 0.0 536.15 0.14 ;
    RECT 535.55 0.0 535.69 0.14 ;
    RECT 534.52 0.0 534.95 0.14 ;
    RECT 533.18 0.0 534.17 0.14 ;
    RECT 531.98 0.0 532.83 0.14 ;
    RECT 531.2 0.0 531.63 0.14 ;
    RECT 529.86 0.0 530.6 0.14 ;
    RECT 529.33 0.0 529.51 0.14 ;
    RECT 528.91 0.0 529.05 0.14 ;
    RECT 527.88 0.0 528.31 0.14 ;
    RECT 526.54 0.0 527.53 0.14 ;
    RECT 525.34 0.0 526.19 0.14 ;
    RECT 524.56 0.0 524.99 0.14 ;
    RECT 523.22 0.0 523.96 0.14 ;
    RECT 522.69 0.0 522.87 0.14 ;
    RECT 522.27 0.0 522.41 0.14 ;
    RECT 521.24 0.0 521.67 0.14 ;
    RECT 519.9 0.0 520.89 0.14 ;
    RECT 518.7 0.0 519.55 0.14 ;
    RECT 517.92 0.0 518.35 0.14 ;
    RECT 516.58 0.0 517.32 0.14 ;
    RECT 516.05 0.0 516.23 0.14 ;
    RECT 515.63 0.0 515.77 0.14 ;
    RECT 514.6 0.0 515.03 0.14 ;
    RECT 513.26 0.0 514.25 0.14 ;
    RECT 512.06 0.0 512.91 0.14 ;
    RECT 511.28 0.0 511.71 0.14 ;
    RECT 509.94 0.0 510.68 0.14 ;
    RECT 509.41 0.0 509.59 0.14 ;
    RECT 508.99 0.0 509.13 0.14 ;
    RECT 507.96 0.0 508.39 0.14 ;
    RECT 506.62 0.0 507.61 0.14 ;
    RECT 505.42 0.0 506.27 0.14 ;
    RECT 504.64 0.0 505.07 0.14 ;
    RECT 503.3 0.0 504.04 0.14 ;
    RECT 502.77 0.0 502.95 0.14 ;
    RECT 502.35 0.0 502.49 0.14 ;
    RECT 501.32 0.0 501.75 0.14 ;
    RECT 499.98 0.0 500.97 0.14 ;
    RECT 498.78 0.0 499.63 0.14 ;
    RECT 498.0 0.0 498.43 0.14 ;
    RECT 496.66 0.0 497.4 0.14 ;
    RECT 496.13 0.0 496.31 0.14 ;
    RECT 495.71 0.0 495.85 0.14 ;
    RECT 494.68 0.0 495.11 0.14 ;
    RECT 493.34 0.0 494.33 0.14 ;
    RECT 492.14 0.0 492.99 0.14 ;
    RECT 491.36 0.0 491.79 0.14 ;
    RECT 490.02 0.0 490.76 0.14 ;
    RECT 489.49 0.0 489.67 0.14 ;
    RECT 489.07 0.0 489.21 0.14 ;
    RECT 488.04 0.0 488.47 0.14 ;
    RECT 486.7 0.0 487.69 0.14 ;
    RECT 485.5 0.0 486.35 0.14 ;
    RECT 484.72 0.0 485.15 0.14 ;
    RECT 483.38 0.0 484.12 0.14 ;
    RECT 482.85 0.0 483.03 0.14 ;
    RECT 482.43 0.0 482.57 0.14 ;
    RECT 481.4 0.0 481.83 0.14 ;
    RECT 480.06 0.0 481.05 0.14 ;
    RECT 478.86 0.0 479.71 0.14 ;
    RECT 478.08 0.0 478.51 0.14 ;
    RECT 476.74 0.0 477.48 0.14 ;
    RECT 476.21 0.0 476.39 0.14 ;
    RECT 475.79 0.0 475.93 0.14 ;
    RECT 474.76 0.0 475.19 0.14 ;
    RECT 473.42 0.0 474.41 0.14 ;
    RECT 472.22 0.0 473.07 0.14 ;
    RECT 471.44 0.0 471.87 0.14 ;
    RECT 470.1 0.0 470.84 0.14 ;
    RECT 469.57 0.0 469.75 0.14 ;
    RECT 469.15 0.0 469.29 0.14 ;
    RECT 468.12 0.0 468.55 0.14 ;
    RECT 466.78 0.0 467.77 0.14 ;
    RECT 465.58 0.0 466.43 0.14 ;
    RECT 464.8 0.0 465.23 0.14 ;
    RECT 463.46 0.0 464.2 0.14 ;
    RECT 462.93 0.0 463.11 0.14 ;
    RECT 462.51 0.0 462.65 0.14 ;
    RECT 461.48 0.0 461.91 0.14 ;
    RECT 460.14 0.0 461.13 0.14 ;
    RECT 458.94 0.0 459.79 0.14 ;
    RECT 458.16 0.0 458.59 0.14 ;
    RECT 456.82 0.0 457.56 0.14 ;
    RECT 456.29 0.0 456.47 0.14 ;
    RECT 455.87 0.0 456.01 0.14 ;
    RECT 454.84 0.0 455.27 0.14 ;
    RECT 453.5 0.0 454.49 0.14 ;
    RECT 452.3 0.0 453.15 0.14 ;
    RECT 451.52 0.0 451.95 0.14 ;
    RECT 450.18 0.0 450.92 0.14 ;
    RECT 449.65 0.0 449.83 0.14 ;
    RECT 449.23 0.0 449.37 0.14 ;
    RECT 448.2 0.0 448.63 0.14 ;
    RECT 446.86 0.0 447.85 0.14 ;
    RECT 445.66 0.0 446.51 0.14 ;
    RECT 444.88 0.0 445.31 0.14 ;
    RECT 443.54 0.0 444.28 0.14 ;
    RECT 443.01 0.0 443.19 0.14 ;
    RECT 442.59 0.0 442.73 0.14 ;
    RECT 441.56 0.0 441.99 0.14 ;
    RECT 440.22 0.0 441.21 0.14 ;
    RECT 439.02 0.0 439.87 0.14 ;
    RECT 428.215 0.0 438.67 0.14 ;
    RECT 427.535 0.0 427.855 0.14 ;
    RECT 424.785 0.0 427.175 0.14 ;
    RECT 419.68 0.0 424.425 0.14 ;
    RECT 418.34 0.0 419.08 0.14 ;
    RECT 417.81 0.0 417.99 0.14 ;
    RECT 417.39 0.0 417.53 0.14 ;
    RECT 416.36 0.0 416.79 0.14 ;
    RECT 415.02 0.0 416.01 0.14 ;
    RECT 413.82 0.0 414.67 0.14 ;
    RECT 413.04 0.0 413.47 0.14 ;
    RECT 411.7 0.0 412.44 0.14 ;
    RECT 411.17 0.0 411.35 0.14 ;
    RECT 410.75 0.0 410.89 0.14 ;
    RECT 409.72 0.0 410.15 0.14 ;
    RECT 408.38 0.0 409.37 0.14 ;
    RECT 407.18 0.0 408.03 0.14 ;
    RECT 406.4 0.0 406.83 0.14 ;
    RECT 405.06 0.0 405.8 0.14 ;
    RECT 404.53 0.0 404.71 0.14 ;
    RECT 404.11 0.0 404.25 0.14 ;
    RECT 403.08 0.0 403.51 0.14 ;
    RECT 401.74 0.0 402.73 0.14 ;
    RECT 400.54 0.0 401.39 0.14 ;
    RECT 399.76 0.0 400.19 0.14 ;
    RECT 398.42 0.0 399.16 0.14 ;
    RECT 397.89 0.0 398.07 0.14 ;
    RECT 397.47 0.0 397.61 0.14 ;
    RECT 396.44 0.0 396.87 0.14 ;
    RECT 395.1 0.0 396.09 0.14 ;
    RECT 393.9 0.0 394.75 0.14 ;
    RECT 393.12 0.0 393.55 0.14 ;
    RECT 391.78 0.0 392.52 0.14 ;
    RECT 391.25 0.0 391.43 0.14 ;
    RECT 390.83 0.0 390.97 0.14 ;
    RECT 389.8 0.0 390.23 0.14 ;
    RECT 388.46 0.0 389.45 0.14 ;
    RECT 387.26 0.0 388.11 0.14 ;
    RECT 386.48 0.0 386.91 0.14 ;
    RECT 385.14 0.0 385.88 0.14 ;
    RECT 384.61 0.0 384.79 0.14 ;
    RECT 384.19 0.0 384.33 0.14 ;
    RECT 383.16 0.0 383.59 0.14 ;
    RECT 381.82 0.0 382.81 0.14 ;
    RECT 380.62 0.0 381.47 0.14 ;
    RECT 379.84 0.0 380.27 0.14 ;
    RECT 378.5 0.0 379.24 0.14 ;
    RECT 377.97 0.0 378.15 0.14 ;
    RECT 377.55 0.0 377.69 0.14 ;
    RECT 376.52 0.0 376.95 0.14 ;
    RECT 375.18 0.0 376.17 0.14 ;
    RECT 373.98 0.0 374.83 0.14 ;
    RECT 373.2 0.0 373.63 0.14 ;
    RECT 371.86 0.0 372.6 0.14 ;
    RECT 371.33 0.0 371.51 0.14 ;
    RECT 370.91 0.0 371.05 0.14 ;
    RECT 369.88 0.0 370.31 0.14 ;
    RECT 368.54 0.0 369.53 0.14 ;
    RECT 367.34 0.0 368.19 0.14 ;
    RECT 366.56 0.0 366.99 0.14 ;
    RECT 365.22 0.0 365.96 0.14 ;
    RECT 364.69 0.0 364.87 0.14 ;
    RECT 364.27 0.0 364.41 0.14 ;
    RECT 363.24 0.0 363.67 0.14 ;
    RECT 361.9 0.0 362.89 0.14 ;
    RECT 360.7 0.0 361.55 0.14 ;
    RECT 359.92 0.0 360.35 0.14 ;
    RECT 358.58 0.0 359.32 0.14 ;
    RECT 358.05 0.0 358.23 0.14 ;
    RECT 357.63 0.0 357.77 0.14 ;
    RECT 356.6 0.0 357.03 0.14 ;
    RECT 355.26 0.0 356.25 0.14 ;
    RECT 354.06 0.0 354.91 0.14 ;
    RECT 353.28 0.0 353.71 0.14 ;
    RECT 351.94 0.0 352.68 0.14 ;
    RECT 351.41 0.0 351.59 0.14 ;
    RECT 350.99 0.0 351.13 0.14 ;
    RECT 349.96 0.0 350.39 0.14 ;
    RECT 348.62 0.0 349.61 0.14 ;
    RECT 347.42 0.0 348.27 0.14 ;
    RECT 346.64 0.0 347.07 0.14 ;
    RECT 345.3 0.0 346.04 0.14 ;
    RECT 344.77 0.0 344.95 0.14 ;
    RECT 344.35 0.0 344.49 0.14 ;
    RECT 343.32 0.0 343.75 0.14 ;
    RECT 341.98 0.0 342.97 0.14 ;
    RECT 340.78 0.0 341.63 0.14 ;
    RECT 340.0 0.0 340.43 0.14 ;
    RECT 338.66 0.0 339.4 0.14 ;
    RECT 338.13 0.0 338.31 0.14 ;
    RECT 337.71 0.0 337.85 0.14 ;
    RECT 336.68 0.0 337.11 0.14 ;
    RECT 335.34 0.0 336.33 0.14 ;
    RECT 334.14 0.0 334.99 0.14 ;
    RECT 333.36 0.0 333.79 0.14 ;
    RECT 332.02 0.0 332.76 0.14 ;
    RECT 331.49 0.0 331.67 0.14 ;
    RECT 331.07 0.0 331.21 0.14 ;
    RECT 330.04 0.0 330.47 0.14 ;
    RECT 328.7 0.0 329.69 0.14 ;
    RECT 327.5 0.0 328.35 0.14 ;
    RECT 326.72 0.0 327.15 0.14 ;
    RECT 325.38 0.0 326.12 0.14 ;
    RECT 324.85 0.0 325.03 0.14 ;
    RECT 324.43 0.0 324.57 0.14 ;
    RECT 323.4 0.0 323.83 0.14 ;
    RECT 322.06 0.0 323.05 0.14 ;
    RECT 320.86 0.0 321.71 0.14 ;
    RECT 320.08 0.0 320.51 0.14 ;
    RECT 318.74 0.0 319.48 0.14 ;
    RECT 318.21 0.0 318.39 0.14 ;
    RECT 317.79 0.0 317.93 0.14 ;
    RECT 316.76 0.0 317.19 0.14 ;
    RECT 315.42 0.0 316.41 0.14 ;
    RECT 314.22 0.0 315.07 0.14 ;
    RECT 313.44 0.0 313.87 0.14 ;
    RECT 312.1 0.0 312.84 0.14 ;
    RECT 311.57 0.0 311.75 0.14 ;
    RECT 311.15 0.0 311.29 0.14 ;
    RECT 310.12 0.0 310.55 0.14 ;
    RECT 308.78 0.0 309.77 0.14 ;
    RECT 307.58 0.0 308.43 0.14 ;
    RECT 306.8 0.0 307.23 0.14 ;
    RECT 305.46 0.0 306.2 0.14 ;
    RECT 304.93 0.0 305.11 0.14 ;
    RECT 304.51 0.0 304.65 0.14 ;
    RECT 303.48 0.0 303.91 0.14 ;
    RECT 302.14 0.0 303.13 0.14 ;
    RECT 300.94 0.0 301.79 0.14 ;
    RECT 300.16 0.0 300.59 0.14 ;
    RECT 298.82 0.0 299.56 0.14 ;
    RECT 298.29 0.0 298.47 0.14 ;
    RECT 297.87 0.0 298.01 0.14 ;
    RECT 296.84 0.0 297.27 0.14 ;
    RECT 295.5 0.0 296.49 0.14 ;
    RECT 294.3 0.0 295.15 0.14 ;
    RECT 293.52 0.0 293.95 0.14 ;
    RECT 292.18 0.0 292.92 0.14 ;
    RECT 291.65 0.0 291.83 0.14 ;
    RECT 291.23 0.0 291.37 0.14 ;
    RECT 290.2 0.0 290.63 0.14 ;
    RECT 288.86 0.0 289.85 0.14 ;
    RECT 287.66 0.0 288.51 0.14 ;
    RECT 285.0 0.0 287.31 0.14 ;
    RECT 283.8 0.0 284.65 0.14 ;
    RECT 282.46 0.0 283.45 0.14 ;
    RECT 281.68 0.0 282.11 0.14 ;
    RECT 280.94 0.0 281.08 0.14 ;
    RECT 280.48 0.0 280.66 0.14 ;
    RECT 279.39 0.0 280.13 0.14 ;
    RECT 278.36 0.0 278.79 0.14 ;
    RECT 277.16 0.0 278.01 0.14 ;
    RECT 275.82 0.0 276.81 0.14 ;
    RECT 275.04 0.0 275.47 0.14 ;
    RECT 274.3 0.0 274.44 0.14 ;
    RECT 273.84 0.0 274.02 0.14 ;
    RECT 272.75 0.0 273.49 0.14 ;
    RECT 271.72 0.0 272.15 0.14 ;
    RECT 270.52 0.0 271.37 0.14 ;
    RECT 269.18 0.0 270.17 0.14 ;
    RECT 268.4 0.0 268.83 0.14 ;
    RECT 267.66 0.0 267.8 0.14 ;
    RECT 267.2 0.0 267.38 0.14 ;
    RECT 266.11 0.0 266.85 0.14 ;
    RECT 265.08 0.0 265.51 0.14 ;
    RECT 263.88 0.0 264.73 0.14 ;
    RECT 262.54 0.0 263.53 0.14 ;
    RECT 261.76 0.0 262.19 0.14 ;
    RECT 261.02 0.0 261.16 0.14 ;
    RECT 260.56 0.0 260.74 0.14 ;
    RECT 259.47 0.0 260.21 0.14 ;
    RECT 258.44 0.0 258.87 0.14 ;
    RECT 257.24 0.0 258.09 0.14 ;
    RECT 255.9 0.0 256.89 0.14 ;
    RECT 255.12 0.0 255.55 0.14 ;
    RECT 254.38 0.0 254.52 0.14 ;
    RECT 253.92 0.0 254.1 0.14 ;
    RECT 252.83 0.0 253.57 0.14 ;
    RECT 251.8 0.0 252.23 0.14 ;
    RECT 250.6 0.0 251.45 0.14 ;
    RECT 249.26 0.0 250.25 0.14 ;
    RECT 248.48 0.0 248.91 0.14 ;
    RECT 247.74 0.0 247.88 0.14 ;
    RECT 247.28 0.0 247.46 0.14 ;
    RECT 246.19 0.0 246.93 0.14 ;
    RECT 245.16 0.0 245.59 0.14 ;
    RECT 243.96 0.0 244.81 0.14 ;
    RECT 242.62 0.0 243.61 0.14 ;
    RECT 241.84 0.0 242.27 0.14 ;
    RECT 241.1 0.0 241.24 0.14 ;
    RECT 240.64 0.0 240.82 0.14 ;
    RECT 239.55 0.0 240.29 0.14 ;
    RECT 238.52 0.0 238.95 0.14 ;
    RECT 237.32 0.0 238.17 0.14 ;
    RECT 235.98 0.0 236.97 0.14 ;
    RECT 235.2 0.0 235.63 0.14 ;
    RECT 234.46 0.0 234.6 0.14 ;
    RECT 234.0 0.0 234.18 0.14 ;
    RECT 232.91 0.0 233.65 0.14 ;
    RECT 231.88 0.0 232.31 0.14 ;
    RECT 230.68 0.0 231.53 0.14 ;
    RECT 229.34 0.0 230.33 0.14 ;
    RECT 228.56 0.0 228.99 0.14 ;
    RECT 227.82 0.0 227.96 0.14 ;
    RECT 227.36 0.0 227.54 0.14 ;
    RECT 226.27 0.0 227.01 0.14 ;
    RECT 225.24 0.0 225.67 0.14 ;
    RECT 224.04 0.0 224.89 0.14 ;
    RECT 222.7 0.0 223.69 0.14 ;
    RECT 221.92 0.0 222.35 0.14 ;
    RECT 221.18 0.0 221.32 0.14 ;
    RECT 220.72 0.0 220.9 0.14 ;
    RECT 219.63 0.0 220.37 0.14 ;
    RECT 218.6 0.0 219.03 0.14 ;
    RECT 217.4 0.0 218.25 0.14 ;
    RECT 216.06 0.0 217.05 0.14 ;
    RECT 215.28 0.0 215.71 0.14 ;
    RECT 214.54 0.0 214.68 0.14 ;
    RECT 214.08 0.0 214.26 0.14 ;
    RECT 212.99 0.0 213.73 0.14 ;
    RECT 211.96 0.0 212.39 0.14 ;
    RECT 210.76 0.0 211.61 0.14 ;
    RECT 209.42 0.0 210.41 0.14 ;
    RECT 208.64 0.0 209.07 0.14 ;
    RECT 207.9 0.0 208.04 0.14 ;
    RECT 207.44 0.0 207.62 0.14 ;
    RECT 206.35 0.0 207.09 0.14 ;
    RECT 205.32 0.0 205.75 0.14 ;
    RECT 204.12 0.0 204.97 0.14 ;
    RECT 202.78 0.0 203.77 0.14 ;
    RECT 202.0 0.0 202.43 0.14 ;
    RECT 201.26 0.0 201.4 0.14 ;
    RECT 200.8 0.0 200.98 0.14 ;
    RECT 199.71 0.0 200.45 0.14 ;
    RECT 198.68 0.0 199.11 0.14 ;
    RECT 197.48 0.0 198.33 0.14 ;
    RECT 196.14 0.0 197.13 0.14 ;
    RECT 195.36 0.0 195.79 0.14 ;
    RECT 194.62 0.0 194.76 0.14 ;
    RECT 194.16 0.0 194.34 0.14 ;
    RECT 193.07 0.0 193.81 0.14 ;
    RECT 192.04 0.0 192.47 0.14 ;
    RECT 190.84 0.0 191.69 0.14 ;
    RECT 189.5 0.0 190.49 0.14 ;
    RECT 188.72 0.0 189.15 0.14 ;
    RECT 187.98 0.0 188.12 0.14 ;
    RECT 187.52 0.0 187.7 0.14 ;
    RECT 186.43 0.0 187.17 0.14 ;
    RECT 185.4 0.0 185.83 0.14 ;
    RECT 184.2 0.0 185.05 0.14 ;
    RECT 182.86 0.0 183.85 0.14 ;
    RECT 182.08 0.0 182.51 0.14 ;
    RECT 181.34 0.0 181.48 0.14 ;
    RECT 180.88 0.0 181.06 0.14 ;
    RECT 179.79 0.0 180.53 0.14 ;
    RECT 178.76 0.0 179.19 0.14 ;
    RECT 177.56 0.0 178.41 0.14 ;
    RECT 176.22 0.0 177.21 0.14 ;
    RECT 175.44 0.0 175.87 0.14 ;
    RECT 174.7 0.0 174.84 0.14 ;
    RECT 174.24 0.0 174.42 0.14 ;
    RECT 173.15 0.0 173.89 0.14 ;
    RECT 172.12 0.0 172.55 0.14 ;
    RECT 170.92 0.0 171.77 0.14 ;
    RECT 169.58 0.0 170.57 0.14 ;
    RECT 168.8 0.0 169.23 0.14 ;
    RECT 168.06 0.0 168.2 0.14 ;
    RECT 167.6 0.0 167.78 0.14 ;
    RECT 166.51 0.0 167.25 0.14 ;
    RECT 165.48 0.0 165.91 0.14 ;
    RECT 164.28 0.0 165.13 0.14 ;
    RECT 162.94 0.0 163.93 0.14 ;
    RECT 162.16 0.0 162.59 0.14 ;
    RECT 161.42 0.0 161.56 0.14 ;
    RECT 160.96 0.0 161.14 0.14 ;
    RECT 159.87 0.0 160.61 0.14 ;
    RECT 158.84 0.0 159.27 0.14 ;
    RECT 157.64 0.0 158.49 0.14 ;
    RECT 156.3 0.0 157.29 0.14 ;
    RECT 155.52 0.0 155.95 0.14 ;
    RECT 154.78 0.0 154.92 0.14 ;
    RECT 154.32 0.0 154.5 0.14 ;
    RECT 153.23 0.0 153.97 0.14 ;
    RECT 147.885 0.0 152.63 0.14 ;
    RECT 145.135 0.0 147.525 0.14 ;
    RECT 144.455 0.0 144.775 0.14 ;
    RECT 133.64 0.0 144.095 0.14 ;
    RECT 132.44 0.0 133.29 0.14 ;
    RECT 131.1 0.0 132.09 0.14 ;
    RECT 130.32 0.0 130.75 0.14 ;
    RECT 129.58 0.0 129.72 0.14 ;
    RECT 129.12 0.0 129.3 0.14 ;
    RECT 128.03 0.0 128.77 0.14 ;
    RECT 127.0 0.0 127.43 0.14 ;
    RECT 125.8 0.0 126.65 0.14 ;
    RECT 124.46 0.0 125.45 0.14 ;
    RECT 123.68 0.0 124.11 0.14 ;
    RECT 122.94 0.0 123.08 0.14 ;
    RECT 122.48 0.0 122.66 0.14 ;
    RECT 121.39 0.0 122.13 0.14 ;
    RECT 120.36 0.0 120.79 0.14 ;
    RECT 119.16 0.0 120.01 0.14 ;
    RECT 117.82 0.0 118.81 0.14 ;
    RECT 117.04 0.0 117.47 0.14 ;
    RECT 116.3 0.0 116.44 0.14 ;
    RECT 115.84 0.0 116.02 0.14 ;
    RECT 114.75 0.0 115.49 0.14 ;
    RECT 113.72 0.0 114.15 0.14 ;
    RECT 112.52 0.0 113.37 0.14 ;
    RECT 111.18 0.0 112.17 0.14 ;
    RECT 110.4 0.0 110.83 0.14 ;
    RECT 109.66 0.0 109.8 0.14 ;
    RECT 109.2 0.0 109.38 0.14 ;
    RECT 108.11 0.0 108.85 0.14 ;
    RECT 107.08 0.0 107.51 0.14 ;
    RECT 105.88 0.0 106.73 0.14 ;
    RECT 104.54 0.0 105.53 0.14 ;
    RECT 103.76 0.0 104.19 0.14 ;
    RECT 103.02 0.0 103.16 0.14 ;
    RECT 102.56 0.0 102.74 0.14 ;
    RECT 101.47 0.0 102.21 0.14 ;
    RECT 100.44 0.0 100.87 0.14 ;
    RECT 99.24 0.0 100.09 0.14 ;
    RECT 97.9 0.0 98.89 0.14 ;
    RECT 97.12 0.0 97.55 0.14 ;
    RECT 96.38 0.0 96.52 0.14 ;
    RECT 95.92 0.0 96.1 0.14 ;
    RECT 94.83 0.0 95.57 0.14 ;
    RECT 93.8 0.0 94.23 0.14 ;
    RECT 92.6 0.0 93.45 0.14 ;
    RECT 91.26 0.0 92.25 0.14 ;
    RECT 90.48 0.0 90.91 0.14 ;
    RECT 89.74 0.0 89.88 0.14 ;
    RECT 89.28 0.0 89.46 0.14 ;
    RECT 88.19 0.0 88.93 0.14 ;
    RECT 87.16 0.0 87.59 0.14 ;
    RECT 85.96 0.0 86.81 0.14 ;
    RECT 84.62 0.0 85.61 0.14 ;
    RECT 83.84 0.0 84.27 0.14 ;
    RECT 83.1 0.0 83.24 0.14 ;
    RECT 82.64 0.0 82.82 0.14 ;
    RECT 81.55 0.0 82.29 0.14 ;
    RECT 80.52 0.0 80.95 0.14 ;
    RECT 79.32 0.0 80.17 0.14 ;
    RECT 77.98 0.0 78.97 0.14 ;
    RECT 77.2 0.0 77.63 0.14 ;
    RECT 76.46 0.0 76.6 0.14 ;
    RECT 76.0 0.0 76.18 0.14 ;
    RECT 74.91 0.0 75.65 0.14 ;
    RECT 73.88 0.0 74.31 0.14 ;
    RECT 72.68 0.0 73.53 0.14 ;
    RECT 71.34 0.0 72.33 0.14 ;
    RECT 70.56 0.0 70.99 0.14 ;
    RECT 69.82 0.0 69.96 0.14 ;
    RECT 69.36 0.0 69.54 0.14 ;
    RECT 68.27 0.0 69.01 0.14 ;
    RECT 67.24 0.0 67.67 0.14 ;
    RECT 66.04 0.0 66.89 0.14 ;
    RECT 64.7 0.0 65.69 0.14 ;
    RECT 63.92 0.0 64.35 0.14 ;
    RECT 63.18 0.0 63.32 0.14 ;
    RECT 62.72 0.0 62.9 0.14 ;
    RECT 61.63 0.0 62.37 0.14 ;
    RECT 60.6 0.0 61.03 0.14 ;
    RECT 59.4 0.0 60.25 0.14 ;
    RECT 58.06 0.0 59.05 0.14 ;
    RECT 57.28 0.0 57.71 0.14 ;
    RECT 56.54 0.0 56.68 0.14 ;
    RECT 56.08 0.0 56.26 0.14 ;
    RECT 54.99 0.0 55.73 0.14 ;
    RECT 53.96 0.0 54.39 0.14 ;
    RECT 52.76 0.0 53.61 0.14 ;
    RECT 51.42 0.0 52.41 0.14 ;
    RECT 50.64 0.0 51.07 0.14 ;
    RECT 49.9 0.0 50.04 0.14 ;
    RECT 49.44 0.0 49.62 0.14 ;
    RECT 48.35 0.0 49.09 0.14 ;
    RECT 47.32 0.0 47.75 0.14 ;
    RECT 46.12 0.0 46.97 0.14 ;
    RECT 44.78 0.0 45.77 0.14 ;
    RECT 44.0 0.0 44.43 0.14 ;
    RECT 43.26 0.0 43.4 0.14 ;
    RECT 42.8 0.0 42.98 0.14 ;
    RECT 41.71 0.0 42.45 0.14 ;
    RECT 40.68 0.0 41.11 0.14 ;
    RECT 39.48 0.0 40.33 0.14 ;
    RECT 38.14 0.0 39.13 0.14 ;
    RECT 37.36 0.0 37.79 0.14 ;
    RECT 36.62 0.0 36.76 0.14 ;
    RECT 36.16 0.0 36.34 0.14 ;
    RECT 35.07 0.0 35.81 0.14 ;
    RECT 34.04 0.0 34.47 0.14 ;
    RECT 32.84 0.0 33.69 0.14 ;
    RECT 31.5 0.0 32.49 0.14 ;
    RECT 30.72 0.0 31.15 0.14 ;
    RECT 29.98 0.0 30.12 0.14 ;
    RECT 29.52 0.0 29.7 0.14 ;
    RECT 28.43 0.0 29.17 0.14 ;
    RECT 27.4 0.0 27.83 0.14 ;
    RECT 26.2 0.0 27.05 0.14 ;
    RECT 24.86 0.0 25.85 0.14 ;
    RECT 24.08 0.0 24.51 0.14 ;
    RECT 23.34 0.0 23.48 0.14 ;
    RECT 22.88 0.0 23.06 0.14 ;
    RECT 21.79 0.0 22.53 0.14 ;
    RECT 20.76 0.0 21.19 0.14 ;
    RECT 19.56 0.0 20.41 0.14 ;
    RECT 18.22 0.0 19.21 0.14 ;
    RECT 17.44 0.0 17.87 0.14 ;
    RECT 16.7 0.0 16.84 0.14 ;
    RECT 16.24 0.0 16.42 0.14 ;
    RECT 15.15 0.0 15.89 0.14 ;
    RECT 14.12 0.0 14.55 0.14 ;
    RECT 12.92 0.0 13.77 0.14 ;
    RECT 11.58 0.0 12.57 0.14 ;
    RECT 10.8 0.0 11.23 0.14 ;
    RECT 10.06 0.0 10.2 0.14 ;
    RECT 9.6 0.0 9.78 0.14 ;
    RECT 8.51 0.0 9.25 0.14 ;
    RECT 7.48 0.0 7.91 0.14 ;
    RECT 6.28 0.0 7.13 0.14 ;
    RECT 4.94 0.0 5.93 0.14 ;
    RECT 4.16 0.0 4.59 0.14 ;
    RECT 3.42 0.0 3.56 0.14 ;
    RECT 2.96 0.0 3.14 0.14 ;
    RECT 1.87 0.0 2.61 0.14 ;
    RECT 0.0 0.0 1.27 0.14 ;
    RECT 571.04 0.14 572.31 145.84 ;
    RECT 569.7 0.14 570.69 145.84 ;
    RECT 568.5 0.14 569.35 145.84 ;
    RECT 567.72 0.14 568.15 145.84 ;
    RECT 566.38 0.14 567.37 145.84 ;
    RECT 565.18 0.14 566.03 145.84 ;
    RECT 564.4 0.14 564.83 145.84 ;
    RECT 563.06 0.14 564.05 145.84 ;
    RECT 561.86 0.14 562.71 145.84 ;
    RECT 561.08 0.14 561.51 145.84 ;
    RECT 559.74 0.14 560.73 145.84 ;
    RECT 558.54 0.14 559.39 145.84 ;
    RECT 557.76 0.14 558.19 145.84 ;
    RECT 556.42 0.14 557.41 145.84 ;
    RECT 555.22 0.14 556.07 145.84 ;
    RECT 554.44 0.14 554.87 145.84 ;
    RECT 553.1 0.14 554.09 145.84 ;
    RECT 551.9 0.14 552.75 145.84 ;
    RECT 551.12 0.14 551.55 145.84 ;
    RECT 549.78 0.14 550.77 145.84 ;
    RECT 548.58 0.14 549.43 145.84 ;
    RECT 547.8 0.14 548.23 145.84 ;
    RECT 546.46 0.14 547.45 145.84 ;
    RECT 545.26 0.14 546.11 145.84 ;
    RECT 544.48 0.14 544.91 145.84 ;
    RECT 543.14 0.14 544.13 145.84 ;
    RECT 541.94 0.14 542.79 145.84 ;
    RECT 541.16 0.14 541.59 145.84 ;
    RECT 539.82 0.14 540.81 145.84 ;
    RECT 538.62 0.14 539.47 145.84 ;
    RECT 537.84 0.14 538.27 145.84 ;
    RECT 536.5 0.14 537.49 145.84 ;
    RECT 535.3 0.14 536.15 145.84 ;
    RECT 534.52 0.14 534.95 145.84 ;
    RECT 533.18 0.14 534.17 145.84 ;
    RECT 531.98 0.14 532.83 145.84 ;
    RECT 531.2 0.14 531.63 145.84 ;
    RECT 529.86 0.14 530.85 145.84 ;
    RECT 528.66 0.14 529.51 145.84 ;
    RECT 527.88 0.14 528.31 145.84 ;
    RECT 526.54 0.14 527.53 145.84 ;
    RECT 525.34 0.14 526.19 145.84 ;
    RECT 524.56 0.14 524.99 145.84 ;
    RECT 523.22 0.14 524.21 145.84 ;
    RECT 522.02 0.14 522.87 145.84 ;
    RECT 521.24 0.14 521.67 145.84 ;
    RECT 519.9 0.14 520.89 145.84 ;
    RECT 518.7 0.14 519.55 145.84 ;
    RECT 517.92 0.14 518.35 145.84 ;
    RECT 516.58 0.14 517.57 145.84 ;
    RECT 515.38 0.14 516.23 145.84 ;
    RECT 514.6 0.14 515.03 145.84 ;
    RECT 513.26 0.14 514.25 145.84 ;
    RECT 512.06 0.14 512.91 145.84 ;
    RECT 511.28 0.14 511.71 145.84 ;
    RECT 509.94 0.14 510.93 145.84 ;
    RECT 508.74 0.14 509.59 145.84 ;
    RECT 507.96 0.14 508.39 145.84 ;
    RECT 506.62 0.14 507.61 145.84 ;
    RECT 505.42 0.14 506.27 145.84 ;
    RECT 504.64 0.14 505.07 145.84 ;
    RECT 503.3 0.14 504.29 145.84 ;
    RECT 502.1 0.14 502.95 145.84 ;
    RECT 501.32 0.14 501.75 145.84 ;
    RECT 499.98 0.14 500.97 145.84 ;
    RECT 498.78 0.14 499.63 145.84 ;
    RECT 498.0 0.14 498.43 145.84 ;
    RECT 496.66 0.14 497.65 145.84 ;
    RECT 495.46 0.14 496.31 145.84 ;
    RECT 494.68 0.14 495.11 145.84 ;
    RECT 493.34 0.14 494.33 145.84 ;
    RECT 492.14 0.14 492.99 145.84 ;
    RECT 491.36 0.14 491.79 145.84 ;
    RECT 490.02 0.14 491.01 145.84 ;
    RECT 488.82 0.14 489.67 145.84 ;
    RECT 488.04 0.14 488.47 145.84 ;
    RECT 486.7 0.14 487.69 145.84 ;
    RECT 485.5 0.14 486.35 145.84 ;
    RECT 484.72 0.14 485.15 145.84 ;
    RECT 483.38 0.14 484.37 145.84 ;
    RECT 482.18 0.14 483.03 145.84 ;
    RECT 481.4 0.14 481.83 145.84 ;
    RECT 480.06 0.14 481.05 145.84 ;
    RECT 478.86 0.14 479.71 145.84 ;
    RECT 478.08 0.14 478.51 145.84 ;
    RECT 476.74 0.14 477.73 145.84 ;
    RECT 475.54 0.14 476.39 145.84 ;
    RECT 474.76 0.14 475.19 145.84 ;
    RECT 473.42 0.14 474.41 145.84 ;
    RECT 472.22 0.14 473.07 145.84 ;
    RECT 471.44 0.14 471.87 145.84 ;
    RECT 470.1 0.14 471.09 145.84 ;
    RECT 468.9 0.14 469.75 145.84 ;
    RECT 468.12 0.14 468.55 145.84 ;
    RECT 466.78 0.14 467.77 145.84 ;
    RECT 465.58 0.14 466.43 145.84 ;
    RECT 464.8 0.14 465.23 145.84 ;
    RECT 463.46 0.14 464.45 145.84 ;
    RECT 462.26 0.14 463.11 145.84 ;
    RECT 461.48 0.14 461.91 145.84 ;
    RECT 460.14 0.14 461.13 145.84 ;
    RECT 458.94 0.14 459.79 145.84 ;
    RECT 458.16 0.14 458.59 145.84 ;
    RECT 456.82 0.14 457.81 145.84 ;
    RECT 455.62 0.14 456.47 145.84 ;
    RECT 454.84 0.14 455.27 145.84 ;
    RECT 453.5 0.14 454.49 145.84 ;
    RECT 452.3 0.14 453.15 145.84 ;
    RECT 451.52 0.14 451.95 145.84 ;
    RECT 450.18 0.14 451.17 145.84 ;
    RECT 448.98 0.14 449.83 145.84 ;
    RECT 448.2 0.14 448.63 145.84 ;
    RECT 446.86 0.14 447.85 145.84 ;
    RECT 445.66 0.14 446.51 145.84 ;
    RECT 444.88 0.14 445.31 145.84 ;
    RECT 443.54 0.14 444.53 145.84 ;
    RECT 442.34 0.14 443.19 145.84 ;
    RECT 441.56 0.14 441.99 145.84 ;
    RECT 440.22 0.14 441.21 145.84 ;
    RECT 439.02 0.14 439.87 145.84 ;
    RECT 428.215 0.14 438.67 145.84 ;
    RECT 427.535 0.14 427.855 145.84 ;
    RECT 424.785 0.14 427.175 145.84 ;
    RECT 419.68 0.14 424.425 145.84 ;
    RECT 418.34 0.14 419.33 145.84 ;
    RECT 417.14 0.14 417.99 145.84 ;
    RECT 416.36 0.14 416.79 145.84 ;
    RECT 415.02 0.14 416.01 145.84 ;
    RECT 413.82 0.14 414.67 145.84 ;
    RECT 413.04 0.14 413.47 145.84 ;
    RECT 411.7 0.14 412.69 145.84 ;
    RECT 410.5 0.14 411.35 145.84 ;
    RECT 409.72 0.14 410.15 145.84 ;
    RECT 408.38 0.14 409.37 145.84 ;
    RECT 407.18 0.14 408.03 145.84 ;
    RECT 406.4 0.14 406.83 145.84 ;
    RECT 405.06 0.14 406.05 145.84 ;
    RECT 403.86 0.14 404.71 145.84 ;
    RECT 403.08 0.14 403.51 145.84 ;
    RECT 401.74 0.14 402.73 145.84 ;
    RECT 400.54 0.14 401.39 145.84 ;
    RECT 399.76 0.14 400.19 145.84 ;
    RECT 398.42 0.14 399.41 145.84 ;
    RECT 397.22 0.14 398.07 145.84 ;
    RECT 396.44 0.14 396.87 145.84 ;
    RECT 395.1 0.14 396.09 145.84 ;
    RECT 393.9 0.14 394.75 145.84 ;
    RECT 393.12 0.14 393.55 145.84 ;
    RECT 391.78 0.14 392.77 145.84 ;
    RECT 390.58 0.14 391.43 145.84 ;
    RECT 389.8 0.14 390.23 145.84 ;
    RECT 388.46 0.14 389.45 145.84 ;
    RECT 387.26 0.14 388.11 145.84 ;
    RECT 386.48 0.14 386.91 145.84 ;
    RECT 385.14 0.14 386.13 145.84 ;
    RECT 383.94 0.14 384.79 145.84 ;
    RECT 383.16 0.14 383.59 145.84 ;
    RECT 381.82 0.14 382.81 145.84 ;
    RECT 380.62 0.14 381.47 145.84 ;
    RECT 379.84 0.14 380.27 145.84 ;
    RECT 378.5 0.14 379.49 145.84 ;
    RECT 377.3 0.14 378.15 145.84 ;
    RECT 376.52 0.14 376.95 145.84 ;
    RECT 375.18 0.14 376.17 145.84 ;
    RECT 373.98 0.14 374.83 145.84 ;
    RECT 373.2 0.14 373.63 145.84 ;
    RECT 371.86 0.14 372.85 145.84 ;
    RECT 370.66 0.14 371.51 145.84 ;
    RECT 369.88 0.14 370.31 145.84 ;
    RECT 368.54 0.14 369.53 145.84 ;
    RECT 367.34 0.14 368.19 145.84 ;
    RECT 366.56 0.14 366.99 145.84 ;
    RECT 365.22 0.14 366.21 145.84 ;
    RECT 364.02 0.14 364.87 145.84 ;
    RECT 363.24 0.14 363.67 145.84 ;
    RECT 361.9 0.14 362.89 145.84 ;
    RECT 360.7 0.14 361.55 145.84 ;
    RECT 359.92 0.14 360.35 145.84 ;
    RECT 358.58 0.14 359.57 145.84 ;
    RECT 357.38 0.14 358.23 145.84 ;
    RECT 356.6 0.14 357.03 145.84 ;
    RECT 355.26 0.14 356.25 145.84 ;
    RECT 354.06 0.14 354.91 145.84 ;
    RECT 353.28 0.14 353.71 145.84 ;
    RECT 351.94 0.14 352.93 145.84 ;
    RECT 350.74 0.14 351.59 145.84 ;
    RECT 349.96 0.14 350.39 145.84 ;
    RECT 348.62 0.14 349.61 145.84 ;
    RECT 347.42 0.14 348.27 145.84 ;
    RECT 346.64 0.14 347.07 145.84 ;
    RECT 345.3 0.14 346.29 145.84 ;
    RECT 344.1 0.14 344.95 145.84 ;
    RECT 343.32 0.14 343.75 145.84 ;
    RECT 341.98 0.14 342.97 145.84 ;
    RECT 340.78 0.14 341.63 145.84 ;
    RECT 340.0 0.14 340.43 145.84 ;
    RECT 338.66 0.14 339.65 145.84 ;
    RECT 337.46 0.14 338.31 145.84 ;
    RECT 336.68 0.14 337.11 145.84 ;
    RECT 335.34 0.14 336.33 145.84 ;
    RECT 334.14 0.14 334.99 145.84 ;
    RECT 333.36 0.14 333.79 145.84 ;
    RECT 332.02 0.14 333.01 145.84 ;
    RECT 330.82 0.14 331.67 145.84 ;
    RECT 330.04 0.14 330.47 145.84 ;
    RECT 328.7 0.14 329.69 145.84 ;
    RECT 327.5 0.14 328.35 145.84 ;
    RECT 326.72 0.14 327.15 145.84 ;
    RECT 325.38 0.14 326.37 145.84 ;
    RECT 324.18 0.14 325.03 145.84 ;
    RECT 323.4 0.14 323.83 145.84 ;
    RECT 322.06 0.14 323.05 145.84 ;
    RECT 320.86 0.14 321.71 145.84 ;
    RECT 320.08 0.14 320.51 145.84 ;
    RECT 318.74 0.14 319.73 145.84 ;
    RECT 317.54 0.14 318.39 145.84 ;
    RECT 316.76 0.14 317.19 145.84 ;
    RECT 315.42 0.14 316.41 145.84 ;
    RECT 314.22 0.14 315.07 145.84 ;
    RECT 313.44 0.14 313.87 145.84 ;
    RECT 312.1 0.14 313.09 145.84 ;
    RECT 310.9 0.14 311.75 145.84 ;
    RECT 310.12 0.14 310.55 145.84 ;
    RECT 308.78 0.14 309.77 145.84 ;
    RECT 307.58 0.14 308.43 145.84 ;
    RECT 306.8 0.14 307.23 145.84 ;
    RECT 305.46 0.14 306.45 145.84 ;
    RECT 304.26 0.14 305.11 145.84 ;
    RECT 303.48 0.14 303.91 145.84 ;
    RECT 302.14 0.14 303.13 145.84 ;
    RECT 300.94 0.14 301.79 145.84 ;
    RECT 300.16 0.14 300.59 145.84 ;
    RECT 298.82 0.14 299.81 145.84 ;
    RECT 297.62 0.14 298.47 145.84 ;
    RECT 296.84 0.14 297.27 145.84 ;
    RECT 295.5 0.14 296.49 145.84 ;
    RECT 294.3 0.14 295.15 145.84 ;
    RECT 293.52 0.14 293.95 145.84 ;
    RECT 292.18 0.14 293.17 145.84 ;
    RECT 290.98 0.14 291.83 145.84 ;
    RECT 290.2 0.14 290.63 145.84 ;
    RECT 288.86 0.14 289.85 145.84 ;
    RECT 287.66 0.14 288.51 145.84 ;
    RECT 285.0 0.14 287.31 145.84 ;
    RECT 283.8 0.14 284.65 145.84 ;
    RECT 282.46 0.14 283.45 145.84 ;
    RECT 281.68 0.14 282.11 145.84 ;
    RECT 280.48 0.14 281.33 145.84 ;
    RECT 279.14 0.14 280.13 145.84 ;
    RECT 278.36 0.14 278.79 145.84 ;
    RECT 277.16 0.14 278.01 145.84 ;
    RECT 275.82 0.14 276.81 145.84 ;
    RECT 275.04 0.14 275.47 145.84 ;
    RECT 273.84 0.14 274.69 145.84 ;
    RECT 272.5 0.14 273.49 145.84 ;
    RECT 271.72 0.14 272.15 145.84 ;
    RECT 270.52 0.14 271.37 145.84 ;
    RECT 269.18 0.14 270.17 145.84 ;
    RECT 268.4 0.14 268.83 145.84 ;
    RECT 267.2 0.14 268.05 145.84 ;
    RECT 265.86 0.14 266.85 145.84 ;
    RECT 265.08 0.14 265.51 145.84 ;
    RECT 263.88 0.14 264.73 145.84 ;
    RECT 262.54 0.14 263.53 145.84 ;
    RECT 261.76 0.14 262.19 145.84 ;
    RECT 260.56 0.14 261.41 145.84 ;
    RECT 259.22 0.14 260.21 145.84 ;
    RECT 258.44 0.14 258.87 145.84 ;
    RECT 257.24 0.14 258.09 145.84 ;
    RECT 255.9 0.14 256.89 145.84 ;
    RECT 255.12 0.14 255.55 145.84 ;
    RECT 253.92 0.14 254.77 145.84 ;
    RECT 252.58 0.14 253.57 145.84 ;
    RECT 251.8 0.14 252.23 145.84 ;
    RECT 250.6 0.14 251.45 145.84 ;
    RECT 249.26 0.14 250.25 145.84 ;
    RECT 248.48 0.14 248.91 145.84 ;
    RECT 247.28 0.14 248.13 145.84 ;
    RECT 245.94 0.14 246.93 145.84 ;
    RECT 245.16 0.14 245.59 145.84 ;
    RECT 243.96 0.14 244.81 145.84 ;
    RECT 242.62 0.14 243.61 145.84 ;
    RECT 241.84 0.14 242.27 145.84 ;
    RECT 240.64 0.14 241.49 145.84 ;
    RECT 239.3 0.14 240.29 145.84 ;
    RECT 238.52 0.14 238.95 145.84 ;
    RECT 237.32 0.14 238.17 145.84 ;
    RECT 235.98 0.14 236.97 145.84 ;
    RECT 235.2 0.14 235.63 145.84 ;
    RECT 234.0 0.14 234.85 145.84 ;
    RECT 232.66 0.14 233.65 145.84 ;
    RECT 231.88 0.14 232.31 145.84 ;
    RECT 230.68 0.14 231.53 145.84 ;
    RECT 229.34 0.14 230.33 145.84 ;
    RECT 228.56 0.14 228.99 145.84 ;
    RECT 227.36 0.14 228.21 145.84 ;
    RECT 226.02 0.14 227.01 145.84 ;
    RECT 225.24 0.14 225.67 145.84 ;
    RECT 224.04 0.14 224.89 145.84 ;
    RECT 222.7 0.14 223.69 145.84 ;
    RECT 221.92 0.14 222.35 145.84 ;
    RECT 220.72 0.14 221.57 145.84 ;
    RECT 219.38 0.14 220.37 145.84 ;
    RECT 218.6 0.14 219.03 145.84 ;
    RECT 217.4 0.14 218.25 145.84 ;
    RECT 216.06 0.14 217.05 145.84 ;
    RECT 215.28 0.14 215.71 145.84 ;
    RECT 214.08 0.14 214.93 145.84 ;
    RECT 212.74 0.14 213.73 145.84 ;
    RECT 211.96 0.14 212.39 145.84 ;
    RECT 210.76 0.14 211.61 145.84 ;
    RECT 209.42 0.14 210.41 145.84 ;
    RECT 208.64 0.14 209.07 145.84 ;
    RECT 207.44 0.14 208.29 145.84 ;
    RECT 206.1 0.14 207.09 145.84 ;
    RECT 205.32 0.14 205.75 145.84 ;
    RECT 204.12 0.14 204.97 145.84 ;
    RECT 202.78 0.14 203.77 145.84 ;
    RECT 202.0 0.14 202.43 145.84 ;
    RECT 200.8 0.14 201.65 145.84 ;
    RECT 199.46 0.14 200.45 145.84 ;
    RECT 198.68 0.14 199.11 145.84 ;
    RECT 197.48 0.14 198.33 145.84 ;
    RECT 196.14 0.14 197.13 145.84 ;
    RECT 195.36 0.14 195.79 145.84 ;
    RECT 194.16 0.14 195.01 145.84 ;
    RECT 192.82 0.14 193.81 145.84 ;
    RECT 192.04 0.14 192.47 145.84 ;
    RECT 190.84 0.14 191.69 145.84 ;
    RECT 189.5 0.14 190.49 145.84 ;
    RECT 188.72 0.14 189.15 145.84 ;
    RECT 187.52 0.14 188.37 145.84 ;
    RECT 186.18 0.14 187.17 145.84 ;
    RECT 185.4 0.14 185.83 145.84 ;
    RECT 184.2 0.14 185.05 145.84 ;
    RECT 182.86 0.14 183.85 145.84 ;
    RECT 182.08 0.14 182.51 145.84 ;
    RECT 180.88 0.14 181.73 145.84 ;
    RECT 179.54 0.14 180.53 145.84 ;
    RECT 178.76 0.14 179.19 145.84 ;
    RECT 177.56 0.14 178.41 145.84 ;
    RECT 176.22 0.14 177.21 145.84 ;
    RECT 175.44 0.14 175.87 145.84 ;
    RECT 174.24 0.14 175.09 145.84 ;
    RECT 172.9 0.14 173.89 145.84 ;
    RECT 172.12 0.14 172.55 145.84 ;
    RECT 170.92 0.14 171.77 145.84 ;
    RECT 169.58 0.14 170.57 145.84 ;
    RECT 168.8 0.14 169.23 145.84 ;
    RECT 167.6 0.14 168.45 145.84 ;
    RECT 166.26 0.14 167.25 145.84 ;
    RECT 165.48 0.14 165.91 145.84 ;
    RECT 164.28 0.14 165.13 145.84 ;
    RECT 162.94 0.14 163.93 145.84 ;
    RECT 162.16 0.14 162.59 145.84 ;
    RECT 160.96 0.14 161.81 145.84 ;
    RECT 159.62 0.14 160.61 145.84 ;
    RECT 158.84 0.14 159.27 145.84 ;
    RECT 157.64 0.14 158.49 145.84 ;
    RECT 156.3 0.14 157.29 145.84 ;
    RECT 155.52 0.14 155.95 145.84 ;
    RECT 154.32 0.14 155.17 145.84 ;
    RECT 152.98 0.14 153.97 145.84 ;
    RECT 147.885 0.14 152.63 145.84 ;
    RECT 145.135 0.14 147.525 145.84 ;
    RECT 144.455 0.14 144.775 145.84 ;
    RECT 133.64 0.14 144.095 145.84 ;
    RECT 132.44 0.14 133.29 145.84 ;
    RECT 131.1 0.14 132.09 145.84 ;
    RECT 130.32 0.14 130.75 145.84 ;
    RECT 129.12 0.14 129.97 145.84 ;
    RECT 127.78 0.14 128.77 145.84 ;
    RECT 127.0 0.14 127.43 145.84 ;
    RECT 125.8 0.14 126.65 145.84 ;
    RECT 124.46 0.14 125.45 145.84 ;
    RECT 123.68 0.14 124.11 145.84 ;
    RECT 122.48 0.14 123.33 145.84 ;
    RECT 121.14 0.14 122.13 145.84 ;
    RECT 120.36 0.14 120.79 145.84 ;
    RECT 119.16 0.14 120.01 145.84 ;
    RECT 117.82 0.14 118.81 145.84 ;
    RECT 117.04 0.14 117.47 145.84 ;
    RECT 115.84 0.14 116.69 145.84 ;
    RECT 114.5 0.14 115.49 145.84 ;
    RECT 113.72 0.14 114.15 145.84 ;
    RECT 112.52 0.14 113.37 145.84 ;
    RECT 111.18 0.14 112.17 145.84 ;
    RECT 110.4 0.14 110.83 145.84 ;
    RECT 109.2 0.14 110.05 145.84 ;
    RECT 107.86 0.14 108.85 145.84 ;
    RECT 107.08 0.14 107.51 145.84 ;
    RECT 105.88 0.14 106.73 145.84 ;
    RECT 104.54 0.14 105.53 145.84 ;
    RECT 103.76 0.14 104.19 145.84 ;
    RECT 102.56 0.14 103.41 145.84 ;
    RECT 101.22 0.14 102.21 145.84 ;
    RECT 100.44 0.14 100.87 145.84 ;
    RECT 99.24 0.14 100.09 145.84 ;
    RECT 97.9 0.14 98.89 145.84 ;
    RECT 97.12 0.14 97.55 145.84 ;
    RECT 95.92 0.14 96.77 145.84 ;
    RECT 94.58 0.14 95.57 145.84 ;
    RECT 93.8 0.14 94.23 145.84 ;
    RECT 92.6 0.14 93.45 145.84 ;
    RECT 91.26 0.14 92.25 145.84 ;
    RECT 90.48 0.14 90.91 145.84 ;
    RECT 89.28 0.14 90.13 145.84 ;
    RECT 87.94 0.14 88.93 145.84 ;
    RECT 87.16 0.14 87.59 145.84 ;
    RECT 85.96 0.14 86.81 145.84 ;
    RECT 84.62 0.14 85.61 145.84 ;
    RECT 83.84 0.14 84.27 145.84 ;
    RECT 82.64 0.14 83.49 145.84 ;
    RECT 81.3 0.14 82.29 145.84 ;
    RECT 80.52 0.14 80.95 145.84 ;
    RECT 79.32 0.14 80.17 145.84 ;
    RECT 77.98 0.14 78.97 145.84 ;
    RECT 77.2 0.14 77.63 145.84 ;
    RECT 76.0 0.14 76.85 145.84 ;
    RECT 74.66 0.14 75.65 145.84 ;
    RECT 73.88 0.14 74.31 145.84 ;
    RECT 72.68 0.14 73.53 145.84 ;
    RECT 71.34 0.14 72.33 145.84 ;
    RECT 70.56 0.14 70.99 145.84 ;
    RECT 69.36 0.14 70.21 145.84 ;
    RECT 68.02 0.14 69.01 145.84 ;
    RECT 67.24 0.14 67.67 145.84 ;
    RECT 66.04 0.14 66.89 145.84 ;
    RECT 64.7 0.14 65.69 145.84 ;
    RECT 63.92 0.14 64.35 145.84 ;
    RECT 62.72 0.14 63.57 145.84 ;
    RECT 61.38 0.14 62.37 145.84 ;
    RECT 60.6 0.14 61.03 145.84 ;
    RECT 59.4 0.14 60.25 145.84 ;
    RECT 58.06 0.14 59.05 145.84 ;
    RECT 57.28 0.14 57.71 145.84 ;
    RECT 56.08 0.14 56.93 145.84 ;
    RECT 54.74 0.14 55.73 145.84 ;
    RECT 53.96 0.14 54.39 145.84 ;
    RECT 52.76 0.14 53.61 145.84 ;
    RECT 51.42 0.14 52.41 145.84 ;
    RECT 50.64 0.14 51.07 145.84 ;
    RECT 49.44 0.14 50.29 145.84 ;
    RECT 48.1 0.14 49.09 145.84 ;
    RECT 47.32 0.14 47.75 145.84 ;
    RECT 46.12 0.14 46.97 145.84 ;
    RECT 44.78 0.14 45.77 145.84 ;
    RECT 44.0 0.14 44.43 145.84 ;
    RECT 42.8 0.14 43.65 145.84 ;
    RECT 41.46 0.14 42.45 145.84 ;
    RECT 40.68 0.14 41.11 145.84 ;
    RECT 39.48 0.14 40.33 145.84 ;
    RECT 38.14 0.14 39.13 145.84 ;
    RECT 37.36 0.14 37.79 145.84 ;
    RECT 36.16 0.14 37.01 145.84 ;
    RECT 34.82 0.14 35.81 145.84 ;
    RECT 34.04 0.14 34.47 145.84 ;
    RECT 32.84 0.14 33.69 145.84 ;
    RECT 31.5 0.14 32.49 145.84 ;
    RECT 30.72 0.14 31.15 145.84 ;
    RECT 29.52 0.14 30.37 145.84 ;
    RECT 28.18 0.14 29.17 145.84 ;
    RECT 27.4 0.14 27.83 145.84 ;
    RECT 26.2 0.14 27.05 145.84 ;
    RECT 24.86 0.14 25.85 145.84 ;
    RECT 24.08 0.14 24.51 145.84 ;
    RECT 22.88 0.14 23.73 145.84 ;
    RECT 21.54 0.14 22.53 145.84 ;
    RECT 20.76 0.14 21.19 145.84 ;
    RECT 19.56 0.14 20.41 145.84 ;
    RECT 18.22 0.14 19.21 145.84 ;
    RECT 17.44 0.14 17.87 145.84 ;
    RECT 16.24 0.14 17.09 145.84 ;
    RECT 14.9 0.14 15.89 145.84 ;
    RECT 14.12 0.14 14.55 145.84 ;
    RECT 12.92 0.14 13.77 145.84 ;
    RECT 11.58 0.14 12.57 145.84 ;
    RECT 10.8 0.14 11.23 145.84 ;
    RECT 9.6 0.14 10.45 145.84 ;
    RECT 8.26 0.14 9.25 145.84 ;
    RECT 7.48 0.14 7.91 145.84 ;
    RECT 6.28 0.14 7.13 145.84 ;
    RECT 4.94 0.14 5.93 145.84 ;
    RECT 4.16 0.14 4.59 145.84 ;
    RECT 2.96 0.14 3.81 145.84 ;
    RECT 1.62 0.14 2.61 145.84 ;
    RECT 0.0 0.14 1.27 145.84 ;
    LAYER OVERLAP ;
    RECT 0.0 0.0 572.31 145.84 ;
    END
  END sram_sp_hde

END LIBRARY

