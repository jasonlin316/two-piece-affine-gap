module shift_register(
    clk,
    data_in,
    data_out
);
input clk;
input  [79:0] data_in;
output [79:0] data_out;

reg [4:0]  d1;
reg [9:0]  d2;
reg [14:0] d3;
reg [19:0] d4;
reg [24:0] d5;
reg [29:0] d6;
reg [34:0] d7;
reg [39:0] d8;
reg [44:0] d9;
reg [49:0] d10;
reg [54:0] d11;
reg [59:0] d12;
reg [64:0] d13;
reg [69:0] d14;
reg [74:0] d15;
reg [79:0] d16;

//assign data_out = {d16[79:75],d15[74:70],d14[69:65],d13[64:60],d12[59:55],d11[54:50],d10[49:45],
//                    d9[44:40],d8[39:35],d7[34:30],d6[29:25],d5[24:20],d4[19:15],d3[14:10],d2[9:5],d1[4:0]};

assign data_out = {d1[4:0],d2[9:5],d3[14:10],d4[19:15],d5[24:20],d6[29:25],d7[34:30],d8[39:35],d9[44:40],d10[49:45],
                    d11[54:50],d12[59:55],d13[64:60],d14[69:65],d15[74:70],d16[79:75]};

always@(posedge clk)
begin
    d2 <= d2 << 5;
    d3 <= d3 << 5;
    d4 <= d4 << 5;
    d5 <= d5 << 5;
    d6 <= d6 << 5;
    d7 <= d7 << 5;
    d8 <= d8 << 5;
    d9 <= d9 << 5;
    d10 <= d10 << 5;
    d11 <= d11 << 5;
    d12 <= d12 << 5;
    d13 <= d13 << 5;
    d14 <= d14 << 5;
    d15 <= d15 << 5;
    d16 <= d16 << 5;

    d1       <= data_in[4:0];
    d2[4:0]  <= data_in[9:5];
    d3[4:0]  <= data_in[14:10];
    d4[4:0]  <= data_in[19:15];
    d5[4:0]  <= data_in[24:20];
    d6[4:0]  <= data_in[29:25];
    d7[4:0]  <= data_in[34:30];
    d8[4:0]  <= data_in[39:35];
    d9[4:0]  <= data_in[44:40];
    d10[4:0] <= data_in[49:45];
    d11[4:0] <= data_in[54:50];
    d12[4:0] <= data_in[59:55];
    d13[4:0] <= data_in[64:60];
    d14[4:0] <= data_in[69:65];
    d15[4:0] <= data_in[74:70];
    d16[4:0] <= data_in[79:75];
end

endmodule