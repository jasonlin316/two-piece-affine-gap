# Confidential Information of ARM, Inc.
# Use subject to ARM license.
# Copyright (c) 2020 ARM, Inc.

# ACI Version r5p0

# Reifier 3.1.1

VERSION 5.6 ;

BUSBITCHARS "[]" ;

#name: High Density Dual Port SRAM RVT-HVT-RVT Compiler|40G 40nm Process, 256 Rows Per Bank, 0.589um^2 Bit Cell
#version: r5p0
#comment: 
#configuration:  -instname "sram_dp_hde" -words 2048 -bits 80 -frequency 100 -mux 4 -pipeline off -write_mask off -wp_size 8 -write_thru off -top_layer "m5-m9" -power_type otc -redundancy off -rcols 2 -rrows 4 -bmux on -ser none -power_gating off -retention on -ema on -atf off -cust_comment "" -bus_notation on -left_bus_delim "[" -right_bus_delim "]" -pwr_gnd_rename "vddpe:VDDPE,vddce:VDDCE,vsse:VSSE" -prefix "" -name_case upper -rows_p_bl 256 -check_instname on -diodes on -drive 6 -dnw off -dpccm on -corners tt_0p90v_0p90v_25c,ss_0p81v_0p81v_m40c,ss_0p81v_0p81v_125c,ffg_0p99v_0p99v_125c,ff_0p99v_0p99v_m40c,ff_0p99v_0p99v_125c
SITE sram_dp_hde
  CLASS  CORE ;
  SIZE 577.18 BY 270.08 ;
  END sram_dp_hde

MACRO sram_dp_hde
  FOREIGN sram_dp_hde 0 0 ;
  SYMMETRY X Y R90 ;
  SITE sram_dp_hde ;
  SIZE 577.18 BY 270.08 ;
  CLASS BLOCK ;
  PIN TQB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 289.35 0.0 289.49 0.39 ;
      LAYER M4 ;
      RECT 289.35 0.0 289.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[40]
  PIN TQB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 287.69 0.0 287.83 0.39 ;
      LAYER M3 ;
      RECT 287.69 0.0 287.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[39]
  PIN TDB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 289.59 0.0 289.73 0.39 ;
      LAYER M4 ;
      RECT 289.59 0.0 289.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[40]
  PIN TDB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 287.45 0.0 287.59 0.39 ;
      LAYER M3 ;
      RECT 287.45 0.0 287.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[39]
  PIN DYB[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 290.14 0.0 290.28 0.39 ;
      LAYER M2 ;
      RECT 290.14 0.0 290.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[40]
  PIN DYB[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 286.9 0.0 287.04 0.39 ;
      LAYER M1 ;
      RECT 286.9 0.0 287.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[39]
  PIN QB[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 290.89 0.0 291.03 0.39 ;
      LAYER M4 ;
      RECT 290.89 0.0 291.03 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[40]
  PIN QB[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 286.15 0.0 286.29 0.39 ;
      LAYER M3 ;
      RECT 286.15 0.0 286.29 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[39]
  PIN DB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 291.88 0.0 292.02 0.39 ;
      LAYER M4 ;
      RECT 291.88 0.0 292.02 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[40]
  PIN DB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 285.16 0.0 285.3 0.39 ;
      LAYER M3 ;
      RECT 285.16 0.0 285.3 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[39]
  PIN DA[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 292.45 0.0 292.59 0.39 ;
      LAYER M4 ;
      RECT 292.45 0.0 292.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[40]
  PIN DA[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 284.59 0.0 284.73 0.39 ;
      LAYER M3 ;
      RECT 284.59 0.0 284.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[39]
  PIN QA[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 293.44 0.0 293.58 0.39 ;
      LAYER M4 ;
      RECT 293.44 0.0 293.58 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[40]
  PIN QA[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 283.6 0.0 283.74 0.39 ;
      LAYER M3 ;
      RECT 283.6 0.0 283.74 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[39]
  PIN AYB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 293.545 0.0 293.685 0.39 ;
      LAYER M2 ;
      RECT 293.545 0.0 293.685 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[0]
  PIN AYA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 283.36 0.0 283.5 0.39 ;
      LAYER M1 ;
      RECT 283.36 0.0 283.5 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[0]
  PIN DYA[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 294.19 0.0 294.33 0.39 ;
      LAYER M2 ;
      RECT 294.19 0.0 294.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[40]
  PIN DYA[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 282.85 0.0 282.99 0.39 ;
      LAYER M1 ;
      RECT 282.85 0.0 282.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[39]
  PIN TDA[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 294.74 0.0 294.88 0.39 ;
      LAYER M4 ;
      RECT 294.74 0.0 294.88 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[40]
  PIN TDA[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 282.3 0.0 282.44 0.39 ;
      LAYER M3 ;
      RECT 282.3 0.0 282.44 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[39]
  PIN TQA[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 294.98 0.0 295.12 0.39 ;
      LAYER M4 ;
      RECT 294.98 0.0 295.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[40]
  PIN TQA[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 282.06 0.0 282.2 0.39 ;
      LAYER M3 ;
      RECT 282.06 0.0 282.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[39]
  PIN TQB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 295.55 0.0 295.69 0.39 ;
      LAYER M4 ;
      RECT 295.55 0.0 295.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[41]
  PIN TQB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 281.49 0.0 281.63 0.39 ;
      LAYER M3 ;
      RECT 281.49 0.0 281.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[38]
  PIN TDB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 295.79 0.0 295.93 0.39 ;
      LAYER M4 ;
      RECT 295.79 0.0 295.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[41]
  PIN TDB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 281.25 0.0 281.39 0.39 ;
      LAYER M3 ;
      RECT 281.25 0.0 281.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[38]
  PIN TAB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 296.04 0.0 296.18 0.39 ;
      LAYER M2 ;
      RECT 296.04 0.0 296.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[0]
  PIN TAA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 281.0 0.0 281.14 0.39 ;
      LAYER M1 ;
      RECT 281.0 0.0 281.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[0]
  PIN DYB[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 296.34 0.0 296.48 0.39 ;
      LAYER M2 ;
      RECT 296.34 0.0 296.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[41]
  PIN DYB[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 280.7 0.0 280.84 0.39 ;
      LAYER M1 ;
      RECT 280.7 0.0 280.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[38]
  PIN QB[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 297.09 0.0 297.23 0.39 ;
      LAYER M4 ;
      RECT 297.09 0.0 297.23 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[41]
  PIN QB[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 279.95 0.0 280.09 0.39 ;
      LAYER M3 ;
      RECT 279.95 0.0 280.09 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[38]
  PIN AB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 297.33 0.0 297.47 0.39 ;
      LAYER M2 ;
      RECT 297.33 0.0 297.47 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[0]
  PIN AA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 279.785 0.0 279.925 0.39 ;
      LAYER M1 ;
      RECT 279.785 0.0 279.925 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[0]
  PIN DB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 298.08 0.0 298.22 0.39 ;
      LAYER M4 ;
      RECT 298.08 0.0 298.22 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[41]
  PIN DB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 278.96 0.0 279.1 0.39 ;
      LAYER M3 ;
      RECT 278.96 0.0 279.1 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[38]
  PIN DA[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 298.65 0.0 298.79 0.39 ;
      LAYER M4 ;
      RECT 298.65 0.0 298.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[41]
  PIN DA[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 278.39 0.0 278.53 0.39 ;
      LAYER M3 ;
      RECT 278.39 0.0 278.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[38]
  PIN AB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 299.49 0.0 299.63 0.39 ;
      LAYER M2 ;
      RECT 299.49 0.0 299.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[1]
  PIN AA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 277.52 0.0 277.66 0.39 ;
      LAYER M1 ;
      RECT 277.52 0.0 277.66 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[1]
  PIN QA[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 299.64 0.0 299.78 0.39 ;
      LAYER M4 ;
      RECT 299.64 0.0 299.78 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[41]
  PIN QA[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 277.4 0.0 277.54 0.39 ;
      LAYER M3 ;
      RECT 277.4 0.0 277.54 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[38]
  PIN DYA[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 300.39 0.0 300.53 0.39 ;
      LAYER M2 ;
      RECT 300.39 0.0 300.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[41]
  PIN DYA[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 276.65 0.0 276.79 0.39 ;
      LAYER M1 ;
      RECT 276.65 0.0 276.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[38]
  PIN TAB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 300.63 0.0 300.77 0.39 ;
      LAYER M2 ;
      RECT 300.63 0.0 300.77 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[1]
  PIN TAA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 276.41 0.0 276.55 0.39 ;
      LAYER M1 ;
      RECT 276.41 0.0 276.55 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[1]
  PIN TDA[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 300.94 0.0 301.08 0.39 ;
      LAYER M4 ;
      RECT 300.94 0.0 301.08 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[41]
  PIN TDA[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 276.1 0.0 276.24 0.39 ;
      LAYER M3 ;
      RECT 276.1 0.0 276.24 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[38]
  PIN TQA[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 301.18 0.0 301.32 0.39 ;
      LAYER M4 ;
      RECT 301.18 0.0 301.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[41]
  PIN TQA[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 275.86 0.0 276.0 0.39 ;
      LAYER M3 ;
      RECT 275.86 0.0 276.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[38]
  PIN TQB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 301.75 0.0 301.89 0.39 ;
      LAYER M4 ;
      RECT 301.75 0.0 301.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[42]
  PIN TQB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 275.29 0.0 275.43 0.39 ;
      LAYER M3 ;
      RECT 275.29 0.0 275.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[37]
  PIN TDB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 301.99 0.0 302.13 0.39 ;
      LAYER M4 ;
      RECT 301.99 0.0 302.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[42]
  PIN TDB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 275.05 0.0 275.19 0.39 ;
      LAYER M3 ;
      RECT 275.05 0.0 275.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[37]
  PIN DYB[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 302.54 0.0 302.68 0.39 ;
      LAYER M2 ;
      RECT 302.54 0.0 302.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[42]
  PIN DYB[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 274.5 0.0 274.64 0.39 ;
      LAYER M1 ;
      RECT 274.5 0.0 274.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[37]
  PIN AYB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 303.13 0.0 303.27 0.39 ;
      LAYER M2 ;
      RECT 303.13 0.0 303.27 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[1]
  PIN AYA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 273.91 0.0 274.05 0.39 ;
      LAYER M1 ;
      RECT 273.91 0.0 274.05 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[1]
  PIN QB[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 303.29 0.0 303.43 0.39 ;
      LAYER M4 ;
      RECT 303.29 0.0 303.43 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[42]
  PIN QB[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 273.75 0.0 273.89 0.39 ;
      LAYER M3 ;
      RECT 273.75 0.0 273.89 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[37]
  PIN DB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 304.28 0.0 304.42 0.39 ;
      LAYER M4 ;
      RECT 304.28 0.0 304.42 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[42]
  PIN DB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 272.76 0.0 272.9 0.39 ;
      LAYER M3 ;
      RECT 272.76 0.0 272.9 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[37]
  PIN DA[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 304.85 0.0 304.99 0.39 ;
      LAYER M4 ;
      RECT 304.85 0.0 304.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[42]
  PIN DA[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 272.19 0.0 272.33 0.39 ;
      LAYER M3 ;
      RECT 272.19 0.0 272.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[37]
  PIN QA[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 305.84 0.0 305.98 0.39 ;
      LAYER M4 ;
      RECT 305.84 0.0 305.98 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[42]
  PIN QA[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 271.2 0.0 271.34 0.39 ;
      LAYER M3 ;
      RECT 271.2 0.0 271.34 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[37]
  PIN DYA[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 306.59 0.0 306.73 0.39 ;
      LAYER M2 ;
      RECT 306.59 0.0 306.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[42]
  PIN COLLDISN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 270.98 0.0 271.12 0.39 ;
      LAYER M1 ;
      RECT 270.98 0.0 271.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END COLLDISN
  PIN TDA[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 307.14 0.0 307.28 0.39 ;
      LAYER M4 ;
      RECT 307.14 0.0 307.28 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[42]
  PIN DYA[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 270.45 0.0 270.59 0.39 ;
      LAYER M1 ;
      RECT 270.45 0.0 270.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[37]
  PIN TQA[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 307.38 0.0 307.52 0.39 ;
      LAYER M4 ;
      RECT 307.38 0.0 307.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[42]
  PIN TDA[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 269.9 0.0 270.04 0.39 ;
      LAYER M3 ;
      RECT 269.9 0.0 270.04 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[37]
  PIN TQB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 307.95 0.0 308.09 0.39 ;
      LAYER M4 ;
      RECT 307.95 0.0 308.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[43]
  PIN TQA[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 269.66 0.0 269.8 0.39 ;
      LAYER M3 ;
      RECT 269.66 0.0 269.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[37]
  PIN TDB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 308.19 0.0 308.33 0.39 ;
      LAYER M4 ;
      RECT 308.19 0.0 308.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[43]
  PIN TQB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 269.09 0.0 269.23 0.39 ;
      LAYER M3 ;
      RECT 269.09 0.0 269.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[36]
  PIN DYB[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 308.74 0.0 308.88 0.39 ;
      LAYER M2 ;
      RECT 308.74 0.0 308.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[43]
  PIN TDB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 268.85 0.0 268.99 0.39 ;
      LAYER M3 ;
      RECT 268.85 0.0 268.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[36]
  PIN QB[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 309.49 0.0 309.63 0.39 ;
      LAYER M4 ;
      RECT 309.49 0.0 309.63 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[43]
  PIN DYB[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 268.3 0.0 268.44 0.39 ;
      LAYER M1 ;
      RECT 268.3 0.0 268.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[36]
  PIN CLKB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 310.465 0.0 310.605 0.39 ;
      LAYER M2 ;
      RECT 310.465 0.0 310.605 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END CLKB
  PIN QB[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 267.55 0.0 267.69 0.39 ;
      LAYER M3 ;
      RECT 267.55 0.0 267.69 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[36]
  PIN DB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 310.48 0.0 310.62 0.39 ;
      LAYER M4 ;
      RECT 310.48 0.0 310.62 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[43]
  PIN DB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 266.56 0.0 266.7 0.39 ;
      LAYER M3 ;
      RECT 266.56 0.0 266.7 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[36]
  PIN DA[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 311.05 0.0 311.19 0.39 ;
      LAYER M4 ;
      RECT 311.05 0.0 311.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[43]
  PIN DA[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.99 0.0 266.13 0.39 ;
      LAYER M3 ;
      RECT 265.99 0.0 266.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[36]
  PIN QA[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 312.04 0.0 312.18 0.39 ;
      LAYER M4 ;
      RECT 312.04 0.0 312.18 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[43]
  PIN QA[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 265.0 0.0 265.14 0.39 ;
      LAYER M3 ;
      RECT 265.0 0.0 265.14 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[36]
  PIN DYA[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 312.79 0.0 312.93 0.39 ;
      LAYER M2 ;
      RECT 312.79 0.0 312.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[43]
  PIN DYA[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 264.25 0.0 264.39 0.39 ;
      LAYER M1 ;
      RECT 264.25 0.0 264.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[36]
  PIN TDA[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 313.34 0.0 313.48 0.39 ;
      LAYER M4 ;
      RECT 313.34 0.0 313.48 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[43]
  PIN TDA[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 263.7 0.0 263.84 0.39 ;
      LAYER M3 ;
      RECT 263.7 0.0 263.84 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[36]
  PIN TQA[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 313.58 0.0 313.72 0.39 ;
      LAYER M4 ;
      RECT 313.58 0.0 313.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[43]
  PIN TQA[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 263.46 0.0 263.6 0.39 ;
      LAYER M3 ;
      RECT 263.46 0.0 263.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[36]
  PIN TQB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 314.15 0.0 314.29 0.39 ;
      LAYER M4 ;
      RECT 314.15 0.0 314.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[44]
  PIN TQB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 262.89 0.0 263.03 0.39 ;
      LAYER M3 ;
      RECT 262.89 0.0 263.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[35]
  PIN TDB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 314.39 0.0 314.53 0.39 ;
      LAYER M4 ;
      RECT 314.39 0.0 314.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[44]
  PIN TDB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 262.65 0.0 262.79 0.39 ;
      LAYER M3 ;
      RECT 262.65 0.0 262.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[35]
  PIN DYB[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 314.94 0.0 315.08 0.39 ;
      LAYER M2 ;
      RECT 314.94 0.0 315.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[44]
  PIN DYB[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 262.1 0.0 262.24 0.39 ;
      LAYER M1 ;
      RECT 262.1 0.0 262.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[35]
  PIN QB[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 315.69 0.0 315.83 0.39 ;
      LAYER M4 ;
      RECT 315.69 0.0 315.83 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[44]
  PIN QB[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 261.35 0.0 261.49 0.39 ;
      LAYER M3 ;
      RECT 261.35 0.0 261.49 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[35]
  PIN DB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 316.68 0.0 316.82 0.39 ;
      LAYER M4 ;
      RECT 316.68 0.0 316.82 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[44]
  PIN DB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 260.36 0.0 260.5 0.39 ;
      LAYER M3 ;
      RECT 260.36 0.0 260.5 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[35]
  PIN DA[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 317.25 0.0 317.39 0.39 ;
      LAYER M4 ;
      RECT 317.25 0.0 317.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[44]
  PIN CLKA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 259.835 0.0 259.975 0.39 ;
      LAYER M1 ;
      RECT 259.835 0.0 259.975 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END CLKA
  PIN QA[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 318.24 0.0 318.38 0.39 ;
      LAYER M4 ;
      RECT 318.24 0.0 318.38 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[44]
  PIN DA[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 259.79 0.0 259.93 0.39 ;
      LAYER M3 ;
      RECT 259.79 0.0 259.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[35]
  PIN DYA[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 318.99 0.0 319.13 0.39 ;
      LAYER M2 ;
      RECT 318.99 0.0 319.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[44]
  PIN QA[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 258.8 0.0 258.94 0.39 ;
      LAYER M3 ;
      RECT 258.8 0.0 258.94 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[35]
  PIN STOVB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 319.255 0.0 319.395 0.39 ;
      LAYER M2 ;
      RECT 319.255 0.0 319.395 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END STOVB
  PIN DYA[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 258.05 0.0 258.19 0.39 ;
      LAYER M1 ;
      RECT 258.05 0.0 258.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[35]
  PIN TDA[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 319.54 0.0 319.68 0.39 ;
      LAYER M4 ;
      RECT 319.54 0.0 319.68 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[44]
  PIN TDA[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 257.5 0.0 257.64 0.39 ;
      LAYER M3 ;
      RECT 257.5 0.0 257.64 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[35]
  PIN TQA[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 319.78 0.0 319.92 0.39 ;
      LAYER M4 ;
      RECT 319.78 0.0 319.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[44]
  PIN TQA[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 257.26 0.0 257.4 0.39 ;
      LAYER M3 ;
      RECT 257.26 0.0 257.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[35]
  PIN EMASB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 319.825 0.0 319.965 0.39 ;
      LAYER M2 ;
      RECT 319.825 0.0 319.965 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMASB
  PIN TQB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 256.69 0.0 256.83 0.39 ;
      LAYER M3 ;
      RECT 256.69 0.0 256.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[34]
  PIN TQB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 320.35 0.0 320.49 0.39 ;
      LAYER M4 ;
      RECT 320.35 0.0 320.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[45]
  PIN TDB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 256.45 0.0 256.59 0.39 ;
      LAYER M3 ;
      RECT 256.45 0.0 256.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[34]
  PIN TDB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 320.59 0.0 320.73 0.39 ;
      LAYER M4 ;
      RECT 320.59 0.0 320.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[45]
  PIN DYB[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 255.9 0.0 256.04 0.39 ;
      LAYER M1 ;
      RECT 255.9 0.0 256.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[34]
  PIN EMAWB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 320.84 0.0 320.98 0.39 ;
      LAYER M2 ;
      RECT 320.84 0.0 320.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAWB[0]
  PIN QB[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 255.15 0.0 255.29 0.39 ;
      LAYER M3 ;
      RECT 255.15 0.0 255.29 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[34]
  PIN DYB[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 321.14 0.0 321.28 0.39 ;
      LAYER M2 ;
      RECT 321.14 0.0 321.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[45]
  PIN DB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 254.16 0.0 254.3 0.39 ;
      LAYER M3 ;
      RECT 254.16 0.0 254.3 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[34]
  PIN EMAWB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 321.79 0.0 321.93 0.39 ;
      LAYER M2 ;
      RECT 321.79 0.0 321.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAWB[1]
  PIN STOVA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 254.09 0.0 254.23 0.39 ;
      LAYER M1 ;
      RECT 254.09 0.0 254.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END STOVA
  PIN QB[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 321.89 0.0 322.03 0.39 ;
      LAYER M4 ;
      RECT 321.89 0.0 322.03 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[45]
  PIN EMASA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 253.83 0.0 253.97 0.39 ;
      LAYER M1 ;
      RECT 253.83 0.0 253.97 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMASA
  PIN DB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 322.88 0.0 323.02 0.39 ;
      LAYER M4 ;
      RECT 322.88 0.0 323.02 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[45]
  PIN DA[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 253.59 0.0 253.73 0.39 ;
      LAYER M3 ;
      RECT 253.59 0.0 253.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[34]
  PIN DA[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 323.45 0.0 323.59 0.39 ;
      LAYER M4 ;
      RECT 323.45 0.0 323.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[45]
  PIN EMAWA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 253.57 0.0 253.71 0.39 ;
      LAYER M1 ;
      RECT 253.57 0.0 253.71 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAWA[0]
  PIN QA[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 324.44 0.0 324.58 0.39 ;
      LAYER M4 ;
      RECT 324.44 0.0 324.58 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[45]
  PIN EMAWA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 252.735 0.0 252.875 0.39 ;
      LAYER M1 ;
      RECT 252.735 0.0 252.875 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAWA[1]
  PIN DYA[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 325.19 0.0 325.33 0.39 ;
      LAYER M2 ;
      RECT 325.19 0.0 325.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[45]
  PIN QA[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 252.6 0.0 252.74 0.39 ;
      LAYER M3 ;
      RECT 252.6 0.0 252.74 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[34]
  PIN TDA[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 325.74 0.0 325.88 0.39 ;
      LAYER M4 ;
      RECT 325.74 0.0 325.88 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[45]
  PIN DYA[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 251.85 0.0 251.99 0.39 ;
      LAYER M1 ;
      RECT 251.85 0.0 251.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[34]
  PIN TQA[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 325.98 0.0 326.12 0.39 ;
      LAYER M4 ;
      RECT 325.98 0.0 326.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[45]
  PIN TDA[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 251.3 0.0 251.44 0.39 ;
      LAYER M3 ;
      RECT 251.3 0.0 251.44 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[34]
  PIN TQB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 326.55 0.0 326.69 0.39 ;
      LAYER M4 ;
      RECT 326.55 0.0 326.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[46]
  PIN TQA[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 251.06 0.0 251.2 0.39 ;
      LAYER M3 ;
      RECT 251.06 0.0 251.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[34]
  PIN TDB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 326.79 0.0 326.93 0.39 ;
      LAYER M4 ;
      RECT 326.79 0.0 326.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[46]
  PIN TQB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 250.49 0.0 250.63 0.39 ;
      LAYER M3 ;
      RECT 250.49 0.0 250.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[33]
  PIN EMAB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 327.045 0.0 327.185 0.39 ;
      LAYER M2 ;
      RECT 327.045 0.0 327.185 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAB[0]
  PIN TDB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 250.25 0.0 250.39 0.39 ;
      LAYER M3 ;
      RECT 250.25 0.0 250.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[33]
  PIN DYB[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 327.34 0.0 327.48 0.39 ;
      LAYER M2 ;
      RECT 327.34 0.0 327.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[46]
  PIN DYB[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 249.7 0.0 249.84 0.39 ;
      LAYER M1 ;
      RECT 249.7 0.0 249.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[33]
  PIN EMAB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 327.92 0.0 328.06 0.39 ;
      LAYER M2 ;
      RECT 327.92 0.0 328.06 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAB[1]
  PIN QB[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 248.95 0.0 249.09 0.39 ;
      LAYER M3 ;
      RECT 248.95 0.0 249.09 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[33]
  PIN QB[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 328.09 0.0 328.23 0.39 ;
      LAYER M4 ;
      RECT 328.09 0.0 328.23 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[46]
  PIN DB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 247.96 0.0 248.1 0.39 ;
      LAYER M3 ;
      RECT 247.96 0.0 248.1 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[33]
  PIN EMAB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 328.27 0.0 328.41 0.39 ;
      LAYER M2 ;
      RECT 328.27 0.0 328.41 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAB[2]
  PIN EMAA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 247.935 0.0 248.075 0.39 ;
      LAYER M1 ;
      RECT 247.935 0.0 248.075 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAA[2]
  PIN DB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 329.08 0.0 329.22 0.39 ;
      LAYER M4 ;
      RECT 329.08 0.0 329.22 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[46]
  PIN EMAA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 247.51 0.0 247.65 0.39 ;
      LAYER M1 ;
      RECT 247.51 0.0 247.65 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAA[1]
  PIN DA[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 329.65 0.0 329.79 0.39 ;
      LAYER M4 ;
      RECT 329.65 0.0 329.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[46]
  PIN DA[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 247.39 0.0 247.53 0.39 ;
      LAYER M3 ;
      RECT 247.39 0.0 247.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[33]
  PIN QA[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 330.64 0.0 330.78 0.39 ;
      LAYER M4 ;
      RECT 330.64 0.0 330.78 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[46]
  PIN EMAA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 246.58 0.0 246.72 0.39 ;
      LAYER M1 ;
      RECT 246.58 0.0 246.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END EMAA[0]
  PIN DYA[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 331.39 0.0 331.53 0.39 ;
      LAYER M2 ;
      RECT 331.39 0.0 331.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[46]
  PIN QA[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 246.4 0.0 246.54 0.39 ;
      LAYER M3 ;
      RECT 246.4 0.0 246.54 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[33]
  PIN TDA[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 331.94 0.0 332.08 0.39 ;
      LAYER M4 ;
      RECT 331.94 0.0 332.08 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[46]
  PIN DYA[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 245.65 0.0 245.79 0.39 ;
      LAYER M1 ;
      RECT 245.65 0.0 245.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[33]
  PIN TQA[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 332.18 0.0 332.32 0.39 ;
      LAYER M4 ;
      RECT 332.18 0.0 332.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[46]
  PIN TDA[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 245.1 0.0 245.24 0.39 ;
      LAYER M3 ;
      RECT 245.1 0.0 245.24 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[33]
  PIN AYB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 332.25 0.0 332.39 0.39 ;
      LAYER M2 ;
      RECT 332.25 0.0 332.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[2]
  PIN TQA[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 244.86 0.0 245.0 0.39 ;
      LAYER M3 ;
      RECT 244.86 0.0 245.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[33]
  PIN TQB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 332.75 0.0 332.89 0.39 ;
      LAYER M4 ;
      RECT 332.75 0.0 332.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[47]
  PIN AYA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 244.79 0.0 244.93 0.39 ;
      LAYER M1 ;
      RECT 244.79 0.0 244.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[2]
  PIN TDB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 332.99 0.0 333.13 0.39 ;
      LAYER M4 ;
      RECT 332.99 0.0 333.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[47]
  PIN TQB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 244.29 0.0 244.43 0.39 ;
      LAYER M3 ;
      RECT 244.29 0.0 244.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[32]
  PIN DYB[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 333.54 0.0 333.68 0.39 ;
      LAYER M2 ;
      RECT 333.54 0.0 333.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[47]
  PIN TDB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 244.05 0.0 244.19 0.39 ;
      LAYER M3 ;
      RECT 244.05 0.0 244.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[32]
  PIN QB[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 334.29 0.0 334.43 0.39 ;
      LAYER M4 ;
      RECT 334.29 0.0 334.43 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[47]
  PIN DYB[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 243.5 0.0 243.64 0.39 ;
      LAYER M1 ;
      RECT 243.5 0.0 243.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[32]
  PIN TAB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 334.445 0.0 334.585 0.39 ;
      LAYER M2 ;
      RECT 334.445 0.0 334.585 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[2]
  PIN QB[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 242.75 0.0 242.89 0.39 ;
      LAYER M3 ;
      RECT 242.75 0.0 242.89 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[32]
  PIN DB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 335.28 0.0 335.42 0.39 ;
      LAYER M4 ;
      RECT 335.28 0.0 335.42 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[47]
  PIN TAA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 242.655 0.0 242.795 0.39 ;
      LAYER M1 ;
      RECT 242.655 0.0 242.795 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[2]
  PIN DA[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 335.85 0.0 335.99 0.39 ;
      LAYER M4 ;
      RECT 335.85 0.0 335.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[47]
  PIN DB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 241.76 0.0 241.9 0.39 ;
      LAYER M3 ;
      RECT 241.76 0.0 241.9 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[32]
  PIN AB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 336.625 0.0 336.765 0.39 ;
      LAYER M2 ;
      RECT 336.625 0.0 336.765 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[2]
  PIN DA[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 241.19 0.0 241.33 0.39 ;
      LAYER M3 ;
      RECT 241.19 0.0 241.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[32]
  PIN QA[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 336.84 0.0 336.98 0.39 ;
      LAYER M4 ;
      RECT 336.84 0.0 336.98 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[47]
  PIN AA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 240.395 0.0 240.535 0.39 ;
      LAYER M1 ;
      RECT 240.395 0.0 240.535 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[2]
  PIN DYA[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 337.59 0.0 337.73 0.39 ;
      LAYER M2 ;
      RECT 337.59 0.0 337.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[47]
  PIN QA[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 240.2 0.0 240.34 0.39 ;
      LAYER M3 ;
      RECT 240.2 0.0 240.34 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[32]
  PIN AB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 337.855 0.0 337.995 0.39 ;
      LAYER M2 ;
      RECT 337.855 0.0 337.995 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[3]
  PIN AA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 240.07 0.0 240.21 0.39 ;
      LAYER M1 ;
      RECT 240.07 0.0 240.21 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[3]
  PIN TDA[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 338.14 0.0 338.28 0.39 ;
      LAYER M4 ;
      RECT 338.14 0.0 338.28 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[47]
  PIN DYA[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 239.45 0.0 239.59 0.39 ;
      LAYER M1 ;
      RECT 239.45 0.0 239.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[32]
  PIN TQA[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 338.38 0.0 338.52 0.39 ;
      LAYER M4 ;
      RECT 338.38 0.0 338.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[47]
  PIN TDA[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 238.9 0.0 239.04 0.39 ;
      LAYER M3 ;
      RECT 238.9 0.0 239.04 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[32]
  PIN TAB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 338.745 0.0 338.885 0.39 ;
      LAYER M2 ;
      RECT 338.745 0.0 338.885 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[3]
  PIN TQA[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 238.66 0.0 238.8 0.39 ;
      LAYER M3 ;
      RECT 238.66 0.0 238.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[32]
  PIN TQB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 338.95 0.0 339.09 0.39 ;
      LAYER M4 ;
      RECT 338.95 0.0 339.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[48]
  PIN TAA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 238.245 0.0 238.385 0.39 ;
      LAYER M1 ;
      RECT 238.245 0.0 238.385 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[3]
  PIN TDB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 339.19 0.0 339.33 0.39 ;
      LAYER M4 ;
      RECT 339.19 0.0 339.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[48]
  PIN TQB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 238.09 0.0 238.23 0.39 ;
      LAYER M3 ;
      RECT 238.09 0.0 238.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[31]
  PIN DYB[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 339.74 0.0 339.88 0.39 ;
      LAYER M2 ;
      RECT 339.74 0.0 339.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[48]
  PIN TDB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 237.85 0.0 237.99 0.39 ;
      LAYER M3 ;
      RECT 237.85 0.0 237.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[31]
  PIN QB[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 340.49 0.0 340.63 0.39 ;
      LAYER M4 ;
      RECT 340.49 0.0 340.63 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[48]
  PIN DYB[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 237.3 0.0 237.44 0.39 ;
      LAYER M1 ;
      RECT 237.3 0.0 237.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[31]
  PIN DB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 341.48 0.0 341.62 0.39 ;
      LAYER M4 ;
      RECT 341.48 0.0 341.62 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[48]
  PIN QB[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 236.55 0.0 236.69 0.39 ;
      LAYER M3 ;
      RECT 236.55 0.0 236.69 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[31]
  PIN AYB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 341.58 0.0 341.72 0.39 ;
      LAYER M2 ;
      RECT 341.58 0.0 341.72 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[3]
  PIN DB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 235.56 0.0 235.7 0.39 ;
      LAYER M3 ;
      RECT 235.56 0.0 235.7 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[31]
  PIN DA[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 342.05 0.0 342.19 0.39 ;
      LAYER M4 ;
      RECT 342.05 0.0 342.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[48]
  PIN AYA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 235.46 0.0 235.6 0.39 ;
      LAYER M1 ;
      RECT 235.46 0.0 235.6 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[3]
  PIN QA[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 343.04 0.0 343.18 0.39 ;
      LAYER M4 ;
      RECT 343.04 0.0 343.18 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[48]
  PIN DA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 234.99 0.0 235.13 0.39 ;
      LAYER M3 ;
      RECT 234.99 0.0 235.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[31]
  PIN DYA[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 343.79 0.0 343.93 0.39 ;
      LAYER M2 ;
      RECT 343.79 0.0 343.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[48]
  PIN QA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 234.0 0.0 234.14 0.39 ;
      LAYER M3 ;
      RECT 234.0 0.0 234.14 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[31]
  PIN TDA[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 344.34 0.0 344.48 0.39 ;
      LAYER M4 ;
      RECT 344.34 0.0 344.48 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[48]
  PIN DYA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 233.25 0.0 233.39 0.39 ;
      LAYER M1 ;
      RECT 233.25 0.0 233.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[31]
  PIN TQA[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 344.58 0.0 344.72 0.39 ;
      LAYER M4 ;
      RECT 344.58 0.0 344.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[48]
  PIN TDA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 232.7 0.0 232.84 0.39 ;
      LAYER M3 ;
      RECT 232.7 0.0 232.84 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[31]
  PIN TQB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 345.15 0.0 345.29 0.39 ;
      LAYER M4 ;
      RECT 345.15 0.0 345.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[49]
  PIN TQA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 232.46 0.0 232.6 0.39 ;
      LAYER M3 ;
      RECT 232.46 0.0 232.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[31]
  PIN TDB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 345.39 0.0 345.53 0.39 ;
      LAYER M4 ;
      RECT 345.39 0.0 345.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[49]
  PIN TQB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 231.89 0.0 232.03 0.39 ;
      LAYER M3 ;
      RECT 231.89 0.0 232.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[30]
  PIN DYB[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 345.94 0.0 346.08 0.39 ;
      LAYER M2 ;
      RECT 345.94 0.0 346.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[49]
  PIN TDB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 231.65 0.0 231.79 0.39 ;
      LAYER M3 ;
      RECT 231.65 0.0 231.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[30]
  PIN QB[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 346.69 0.0 346.83 0.39 ;
      LAYER M4 ;
      RECT 346.69 0.0 346.83 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[49]
  PIN DYB[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 231.1 0.0 231.24 0.39 ;
      LAYER M1 ;
      RECT 231.1 0.0 231.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[30]
  PIN DB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 347.68 0.0 347.82 0.39 ;
      LAYER M4 ;
      RECT 347.68 0.0 347.82 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[49]
  PIN QB[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 230.35 0.0 230.49 0.39 ;
      LAYER M3 ;
      RECT 230.35 0.0 230.49 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[30]
  PIN DA[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 348.25 0.0 348.39 0.39 ;
      LAYER M4 ;
      RECT 348.25 0.0 348.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[49]
  PIN DB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 229.36 0.0 229.5 0.39 ;
      LAYER M3 ;
      RECT 229.36 0.0 229.5 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[30]
  PIN QA[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 349.24 0.0 349.38 0.39 ;
      LAYER M4 ;
      RECT 349.24 0.0 349.38 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[49]
  PIN DA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 228.79 0.0 228.93 0.39 ;
      LAYER M3 ;
      RECT 228.79 0.0 228.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[30]
  PIN DYA[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 349.99 0.0 350.13 0.39 ;
      LAYER M2 ;
      RECT 349.99 0.0 350.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[49]
  PIN QA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 227.8 0.0 227.94 0.39 ;
      LAYER M3 ;
      RECT 227.8 0.0 227.94 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[30]
  PIN TDA[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 350.54 0.0 350.68 0.39 ;
      LAYER M4 ;
      RECT 350.54 0.0 350.68 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[49]
  PIN DYA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 227.05 0.0 227.19 0.39 ;
      LAYER M1 ;
      RECT 227.05 0.0 227.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[30]
  PIN TQA[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 350.78 0.0 350.92 0.39 ;
      LAYER M4 ;
      RECT 350.78 0.0 350.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[49]
  PIN TDA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 226.5 0.0 226.64 0.39 ;
      LAYER M3 ;
      RECT 226.5 0.0 226.64 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[30]
  PIN AYB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 351.345 0.0 351.485 0.39 ;
      LAYER M2 ;
      RECT 351.345 0.0 351.485 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[4]
  PIN TQA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 226.26 0.0 226.4 0.39 ;
      LAYER M3 ;
      RECT 226.26 0.0 226.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[30]
  PIN TQB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 351.35 0.0 351.49 0.39 ;
      LAYER M4 ;
      RECT 351.35 0.0 351.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[50]
  PIN AYA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 225.77 0.0 225.91 0.39 ;
      LAYER M1 ;
      RECT 225.77 0.0 225.91 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[4]
  PIN TDB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 351.59 0.0 351.73 0.39 ;
      LAYER M4 ;
      RECT 351.59 0.0 351.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[50]
  PIN TQB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 225.69 0.0 225.83 0.39 ;
      LAYER M3 ;
      RECT 225.69 0.0 225.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[29]
  PIN DYB[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 352.14 0.0 352.28 0.39 ;
      LAYER M2 ;
      RECT 352.14 0.0 352.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[50]
  PIN TDB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 225.45 0.0 225.59 0.39 ;
      LAYER M3 ;
      RECT 225.45 0.0 225.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[29]
  PIN QB[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 352.89 0.0 353.03 0.39 ;
      LAYER M4 ;
      RECT 352.89 0.0 353.03 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[50]
  PIN DYB[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 224.9 0.0 225.04 0.39 ;
      LAYER M1 ;
      RECT 224.9 0.0 225.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[29]
  PIN DB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 353.88 0.0 354.02 0.39 ;
      LAYER M4 ;
      RECT 353.88 0.0 354.02 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[50]
  PIN QB[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 224.15 0.0 224.29 0.39 ;
      LAYER M3 ;
      RECT 224.15 0.0 224.29 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[29]
  PIN TAB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 354.32 0.0 354.46 0.39 ;
      LAYER M2 ;
      RECT 354.32 0.0 354.46 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[4]
  PIN DB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 223.16 0.0 223.3 0.39 ;
      LAYER M3 ;
      RECT 223.16 0.0 223.3 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[29]
  PIN DA[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 354.45 0.0 354.59 0.39 ;
      LAYER M4 ;
      RECT 354.45 0.0 354.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[50]
  PIN TAA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 222.715 0.0 222.855 0.39 ;
      LAYER M1 ;
      RECT 222.715 0.0 222.855 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[4]
  PIN QA[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 355.44 0.0 355.58 0.39 ;
      LAYER M4 ;
      RECT 355.44 0.0 355.58 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[50]
  PIN DA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 222.59 0.0 222.73 0.39 ;
      LAYER M3 ;
      RECT 222.59 0.0 222.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[29]
  PIN AB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 355.585 0.0 355.725 0.39 ;
      LAYER M2 ;
      RECT 355.585 0.0 355.725 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[4]
  PIN QA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 221.6 0.0 221.74 0.39 ;
      LAYER M3 ;
      RECT 221.6 0.0 221.74 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[29]
  PIN DYA[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 356.19 0.0 356.33 0.39 ;
      LAYER M2 ;
      RECT 356.19 0.0 356.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[50]
  PIN DYA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 220.85 0.0 220.99 0.39 ;
      LAYER M1 ;
      RECT 220.85 0.0 220.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[29]
  PIN AB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 356.515 0.0 356.655 0.39 ;
      LAYER M2 ;
      RECT 356.515 0.0 356.655 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[5]
  PIN AA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 220.59 0.0 220.73 0.39 ;
      LAYER M1 ;
      RECT 220.59 0.0 220.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[4]
  PIN TDA[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 356.74 0.0 356.88 0.39 ;
      LAYER M4 ;
      RECT 356.74 0.0 356.88 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[50]
  PIN TDA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 220.3 0.0 220.44 0.39 ;
      LAYER M3 ;
      RECT 220.3 0.0 220.44 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[29]
  PIN TQA[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 356.98 0.0 357.12 0.39 ;
      LAYER M4 ;
      RECT 356.98 0.0 357.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[50]
  PIN TQA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 220.06 0.0 220.2 0.39 ;
      LAYER M3 ;
      RECT 220.06 0.0 220.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[29]
  PIN RET1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 357.13 0.0 357.27 0.39 ;
      LAYER M2 ;
      RECT 357.13 0.0 357.27 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END RET1N
  PIN AA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 219.95 0.0 220.09 0.39 ;
      LAYER M1 ;
      RECT 219.95 0.0 220.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[5]
  PIN TQB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 357.55 0.0 357.69 0.39 ;
      LAYER M4 ;
      RECT 357.55 0.0 357.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[51]
  PIN TQB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 219.49 0.0 219.63 0.39 ;
      LAYER M3 ;
      RECT 219.49 0.0 219.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[28]
  PIN TDB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 357.79 0.0 357.93 0.39 ;
      LAYER M4 ;
      RECT 357.79 0.0 357.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[51]
  PIN TDB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 219.25 0.0 219.39 0.39 ;
      LAYER M3 ;
      RECT 219.25 0.0 219.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[28]
  PIN DYB[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 358.34 0.0 358.48 0.39 ;
      LAYER M2 ;
      RECT 358.34 0.0 358.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[51]
  PIN DYB[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 218.7 0.0 218.84 0.39 ;
      LAYER M1 ;
      RECT 218.7 0.0 218.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[28]
  PIN TAB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 359.01 0.0 359.15 0.39 ;
      LAYER M2 ;
      RECT 359.01 0.0 359.15 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[5]
  PIN TAA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 218.03 0.0 218.17 0.39 ;
      LAYER M1 ;
      RECT 218.03 0.0 218.17 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[5]
  PIN QB[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 359.09 0.0 359.23 0.39 ;
      LAYER M4 ;
      RECT 359.09 0.0 359.23 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[51]
  PIN QB[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 217.95 0.0 218.09 0.39 ;
      LAYER M3 ;
      RECT 217.95 0.0 218.09 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[28]
  PIN DB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 360.08 0.0 360.22 0.39 ;
      LAYER M4 ;
      RECT 360.08 0.0 360.22 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[51]
  PIN DB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 216.96 0.0 217.1 0.39 ;
      LAYER M3 ;
      RECT 216.96 0.0 217.1 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[28]
  PIN DA[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 360.65 0.0 360.79 0.39 ;
      LAYER M4 ;
      RECT 360.65 0.0 360.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[51]
  PIN DA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 216.39 0.0 216.53 0.39 ;
      LAYER M3 ;
      RECT 216.39 0.0 216.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[28]
  PIN AYB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 361.53 0.0 361.67 0.39 ;
      LAYER M2 ;
      RECT 361.53 0.0 361.67 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[5]
  PIN AYA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 215.51 0.0 215.65 0.39 ;
      LAYER M1 ;
      RECT 215.51 0.0 215.65 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[5]
  PIN QA[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 361.64 0.0 361.78 0.39 ;
      LAYER M4 ;
      RECT 361.64 0.0 361.78 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[51]
  PIN QA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 215.4 0.0 215.54 0.39 ;
      LAYER M3 ;
      RECT 215.4 0.0 215.54 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[28]
  PIN DYA[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 362.39 0.0 362.53 0.39 ;
      LAYER M2 ;
      RECT 362.39 0.0 362.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[51]
  PIN DYA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 214.65 0.0 214.79 0.39 ;
      LAYER M1 ;
      RECT 214.65 0.0 214.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[28]
  PIN TDA[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 362.94 0.0 363.08 0.39 ;
      LAYER M4 ;
      RECT 362.94 0.0 363.08 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[51]
  PIN TDA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 214.1 0.0 214.24 0.39 ;
      LAYER M3 ;
      RECT 214.1 0.0 214.24 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[28]
  PIN TQA[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 363.18 0.0 363.32 0.39 ;
      LAYER M4 ;
      RECT 363.18 0.0 363.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[51]
  PIN TQA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 213.86 0.0 214.0 0.39 ;
      LAYER M3 ;
      RECT 213.86 0.0 214.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[28]
  PIN TQB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 363.75 0.0 363.89 0.39 ;
      LAYER M4 ;
      RECT 363.75 0.0 363.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[52]
  PIN TQB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 213.29 0.0 213.43 0.39 ;
      LAYER M3 ;
      RECT 213.29 0.0 213.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[27]
  PIN TDB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 363.99 0.0 364.13 0.39 ;
      LAYER M4 ;
      RECT 363.99 0.0 364.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[52]
  PIN TDB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 213.05 0.0 213.19 0.39 ;
      LAYER M3 ;
      RECT 213.05 0.0 213.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[27]
  PIN DYB[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 364.54 0.0 364.68 0.39 ;
      LAYER M2 ;
      RECT 364.54 0.0 364.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[52]
  PIN DYB[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 212.5 0.0 212.64 0.39 ;
      LAYER M1 ;
      RECT 212.5 0.0 212.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[27]
  PIN QB[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 365.29 0.0 365.43 0.39 ;
      LAYER M4 ;
      RECT 365.29 0.0 365.43 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[52]
  PIN QB[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 211.75 0.0 211.89 0.39 ;
      LAYER M3 ;
      RECT 211.75 0.0 211.89 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[27]
  PIN DB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 366.28 0.0 366.42 0.39 ;
      LAYER M4 ;
      RECT 366.28 0.0 366.42 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[52]
  PIN DB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 210.76 0.0 210.9 0.39 ;
      LAYER M3 ;
      RECT 210.76 0.0 210.9 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[27]
  PIN DA[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 366.85 0.0 366.99 0.39 ;
      LAYER M4 ;
      RECT 366.85 0.0 366.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[52]
  PIN DA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 210.19 0.0 210.33 0.39 ;
      LAYER M3 ;
      RECT 210.19 0.0 210.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[27]
  PIN QA[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 367.84 0.0 367.98 0.39 ;
      LAYER M4 ;
      RECT 367.84 0.0 367.98 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[52]
  PIN QA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 209.2 0.0 209.34 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[27]
  PIN DYA[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 368.59 0.0 368.73 0.39 ;
      LAYER M2 ;
      RECT 368.59 0.0 368.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[52]
  PIN DYA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 208.45 0.0 208.59 0.39 ;
      LAYER M1 ;
      RECT 208.45 0.0 208.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[27]
  PIN TDA[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 369.14 0.0 369.28 0.39 ;
      LAYER M4 ;
      RECT 369.14 0.0 369.28 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[52]
  PIN TDA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 207.9 0.0 208.04 0.39 ;
      LAYER M3 ;
      RECT 207.9 0.0 208.04 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[27]
  PIN TQA[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 369.38 0.0 369.52 0.39 ;
      LAYER M4 ;
      RECT 369.38 0.0 369.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[52]
  PIN TQA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 207.66 0.0 207.8 0.39 ;
      LAYER M3 ;
      RECT 207.66 0.0 207.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[27]
  PIN TQB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 369.95 0.0 370.09 0.39 ;
      LAYER M4 ;
      RECT 369.95 0.0 370.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[53]
  PIN TQB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 207.09 0.0 207.23 0.39 ;
      LAYER M3 ;
      RECT 207.09 0.0 207.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[26]
  PIN TDB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 370.19 0.0 370.33 0.39 ;
      LAYER M4 ;
      RECT 370.19 0.0 370.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[53]
  PIN TDB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 206.85 0.0 206.99 0.39 ;
      LAYER M3 ;
      RECT 206.85 0.0 206.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[26]
  PIN AYB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 370.455 0.0 370.595 0.39 ;
      LAYER M2 ;
      RECT 370.455 0.0 370.595 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[6]
  PIN AYA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 206.575 0.0 206.715 0.39 ;
      LAYER M1 ;
      RECT 206.575 0.0 206.715 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[6]
  PIN DYB[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 370.74 0.0 370.88 0.39 ;
      LAYER M2 ;
      RECT 370.74 0.0 370.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[53]
  PIN DYB[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 206.3 0.0 206.44 0.39 ;
      LAYER M1 ;
      RECT 206.3 0.0 206.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[26]
  PIN QB[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 371.49 0.0 371.63 0.39 ;
      LAYER M4 ;
      RECT 371.49 0.0 371.63 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[53]
  PIN QB[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 205.55 0.0 205.69 0.39 ;
      LAYER M3 ;
      RECT 205.55 0.0 205.69 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[26]
  PIN DB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 372.48 0.0 372.62 0.39 ;
      LAYER M4 ;
      RECT 372.48 0.0 372.62 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[53]
  PIN DB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 204.56 0.0 204.7 0.39 ;
      LAYER M3 ;
      RECT 204.56 0.0 204.7 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[26]
  PIN DA[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 373.05 0.0 373.19 0.39 ;
      LAYER M4 ;
      RECT 373.05 0.0 373.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[53]
  PIN DA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 203.99 0.0 204.13 0.39 ;
      LAYER M3 ;
      RECT 203.99 0.0 204.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[26]
  PIN TAB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 373.98 0.0 374.12 0.39 ;
      LAYER M2 ;
      RECT 373.98 0.0 374.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[6]
  PIN TAA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 203.095 0.0 203.235 0.39 ;
      LAYER M1 ;
      RECT 203.095 0.0 203.235 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[6]
  PIN QA[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 374.04 0.0 374.18 0.39 ;
      LAYER M4 ;
      RECT 374.04 0.0 374.18 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[53]
  PIN QA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 203.0 0.0 203.14 0.39 ;
      LAYER M3 ;
      RECT 203.0 0.0 203.14 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[26]
  PIN DYA[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 374.79 0.0 374.93 0.39 ;
      LAYER M2 ;
      RECT 374.79 0.0 374.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[53]
  PIN DYA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 202.25 0.0 202.39 0.39 ;
      LAYER M1 ;
      RECT 202.25 0.0 202.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[26]
  PIN TDA[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 375.34 0.0 375.48 0.39 ;
      LAYER M4 ;
      RECT 375.34 0.0 375.48 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[53]
  PIN TDA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 201.7 0.0 201.84 0.39 ;
      LAYER M3 ;
      RECT 201.7 0.0 201.84 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[26]
  PIN AB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 375.575 0.0 375.715 0.39 ;
      LAYER M2 ;
      RECT 375.575 0.0 375.715 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[6]
  PIN TQA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 201.46 0.0 201.6 0.39 ;
      LAYER M3 ;
      RECT 201.46 0.0 201.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[26]
  PIN TQA[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 375.58 0.0 375.72 0.39 ;
      LAYER M4 ;
      RECT 375.58 0.0 375.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[53]
  PIN AA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 201.405 0.0 201.545 0.39 ;
      LAYER M1 ;
      RECT 201.405 0.0 201.545 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[6]
  PIN AB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 375.835 0.0 375.975 0.39 ;
      LAYER M2 ;
      RECT 375.835 0.0 375.975 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[7]
  PIN AA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 201.065 0.0 201.205 0.39 ;
      LAYER M1 ;
      RECT 201.065 0.0 201.205 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[7]
  PIN AB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 376.095 0.0 376.235 0.39 ;
      LAYER M2 ;
      RECT 376.095 0.0 376.235 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[8]
  PIN TQB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 200.89 0.0 201.03 0.39 ;
      LAYER M3 ;
      RECT 200.89 0.0 201.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[25]
  PIN TQB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 376.15 0.0 376.29 0.39 ;
      LAYER M4 ;
      RECT 376.15 0.0 376.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[54]
  PIN TDB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 200.65 0.0 200.79 0.39 ;
      LAYER M3 ;
      RECT 200.65 0.0 200.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[25]
  PIN TDB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 376.39 0.0 376.53 0.39 ;
      LAYER M4 ;
      RECT 376.39 0.0 376.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[54]
  PIN AA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 200.375 0.0 200.515 0.39 ;
      LAYER M1 ;
      RECT 200.375 0.0 200.515 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[8]
  PIN DYB[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 376.94 0.0 377.08 0.39 ;
      LAYER M2 ;
      RECT 376.94 0.0 377.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[54]
  PIN DYB[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 200.1 0.0 200.24 0.39 ;
      LAYER M1 ;
      RECT 200.1 0.0 200.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[25]
  PIN QB[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 377.69 0.0 377.83 0.39 ;
      LAYER M4 ;
      RECT 377.69 0.0 377.83 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[54]
  PIN QB[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 199.35 0.0 199.49 0.39 ;
      LAYER M3 ;
      RECT 199.35 0.0 199.49 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[25]
  PIN TAB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 377.78 0.0 377.92 0.39 ;
      LAYER M2 ;
      RECT 377.78 0.0 377.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[8]
  PIN TAA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 199.26 0.0 199.4 0.39 ;
      LAYER M1 ;
      RECT 199.26 0.0 199.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[8]
  PIN DB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 378.68 0.0 378.82 0.39 ;
      LAYER M4 ;
      RECT 378.68 0.0 378.82 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[54]
  PIN DB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 198.36 0.0 198.5 0.39 ;
      LAYER M3 ;
      RECT 198.36 0.0 198.5 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[25]
  PIN TAB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 378.71 0.0 378.85 0.39 ;
      LAYER M2 ;
      RECT 378.71 0.0 378.85 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[7]
  PIN TAA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 198.195 0.0 198.335 0.39 ;
      LAYER M1 ;
      RECT 198.195 0.0 198.335 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[7]
  PIN DA[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 379.25 0.0 379.39 0.39 ;
      LAYER M4 ;
      RECT 379.25 0.0 379.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[54]
  PIN DA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 197.79 0.0 197.93 0.39 ;
      LAYER M3 ;
      RECT 197.79 0.0 197.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[25]
  PIN QA[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 380.24 0.0 380.38 0.39 ;
      LAYER M4 ;
      RECT 380.24 0.0 380.38 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[54]
  PIN QA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 196.8 0.0 196.94 0.39 ;
      LAYER M3 ;
      RECT 196.8 0.0 196.94 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[25]
  PIN AYB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 380.45 0.0 380.59 0.39 ;
      LAYER M2 ;
      RECT 380.45 0.0 380.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[7]
  PIN AYA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 196.6 0.0 196.74 0.39 ;
      LAYER M1 ;
      RECT 196.6 0.0 196.74 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[7]
  PIN DYA[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 380.99 0.0 381.13 0.39 ;
      LAYER M2 ;
      RECT 380.99 0.0 381.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[54]
  PIN DYA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 196.05 0.0 196.19 0.39 ;
      LAYER M1 ;
      RECT 196.05 0.0 196.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[25]
  PIN AYB[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 381.265 0.0 381.405 0.39 ;
      LAYER M2 ;
      RECT 381.265 0.0 381.405 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[8]
  PIN AYA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 195.79 0.0 195.93 0.39 ;
      LAYER M1 ;
      RECT 195.79 0.0 195.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[8]
  PIN TDA[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 381.54 0.0 381.68 0.39 ;
      LAYER M4 ;
      RECT 381.54 0.0 381.68 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[54]
  PIN TDA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 195.5 0.0 195.64 0.39 ;
      LAYER M3 ;
      RECT 195.5 0.0 195.64 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[25]
  PIN TQA[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 381.78 0.0 381.92 0.39 ;
      LAYER M4 ;
      RECT 381.78 0.0 381.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[54]
  PIN TQA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 195.26 0.0 195.4 0.39 ;
      LAYER M3 ;
      RECT 195.26 0.0 195.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[25]
  PIN TENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 382.32 0.0 382.46 0.39 ;
      LAYER M2 ;
      RECT 382.32 0.0 382.46 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TENB
  PIN TENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 194.72 0.0 194.86 0.39 ;
      LAYER M1 ;
      RECT 194.72 0.0 194.86 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TENA
  PIN TQB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 382.35 0.0 382.49 0.39 ;
      LAYER M4 ;
      RECT 382.35 0.0 382.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[55]
  PIN TQB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 194.69 0.0 194.83 0.39 ;
      LAYER M3 ;
      RECT 194.69 0.0 194.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[24]
  PIN TDB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 382.59 0.0 382.73 0.39 ;
      LAYER M4 ;
      RECT 382.59 0.0 382.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[55]
  PIN TDB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 194.45 0.0 194.59 0.39 ;
      LAYER M3 ;
      RECT 194.45 0.0 194.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[24]
  PIN DYB[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 383.14 0.0 383.28 0.39 ;
      LAYER M2 ;
      RECT 383.14 0.0 383.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[55]
  PIN DYB[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 193.9 0.0 194.04 0.39 ;
      LAYER M1 ;
      RECT 193.9 0.0 194.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[24]
  PIN QB[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 383.89 0.0 384.03 0.39 ;
      LAYER M4 ;
      RECT 383.89 0.0 384.03 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[55]
  PIN QB[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 193.15 0.0 193.29 0.39 ;
      LAYER M3 ;
      RECT 193.15 0.0 193.29 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[24]
  PIN DB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 384.88 0.0 385.02 0.39 ;
      LAYER M4 ;
      RECT 384.88 0.0 385.02 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[55]
  PIN DB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 192.16 0.0 192.3 0.39 ;
      LAYER M3 ;
      RECT 192.16 0.0 192.3 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[24]
  PIN BENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 385.4 0.0 385.54 0.39 ;
      LAYER M2 ;
      RECT 385.4 0.0 385.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END BENB
  PIN BENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 191.64 0.0 191.78 0.39 ;
      LAYER M1 ;
      RECT 191.64 0.0 191.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END BENA
  PIN DA[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 385.45 0.0 385.59 0.39 ;
      LAYER M4 ;
      RECT 385.45 0.0 385.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[55]
  PIN DA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 191.59 0.0 191.73 0.39 ;
      LAYER M3 ;
      RECT 191.59 0.0 191.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[24]
  PIN QA[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 386.44 0.0 386.58 0.39 ;
      LAYER M4 ;
      RECT 386.44 0.0 386.58 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[55]
  PIN QA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 190.6 0.0 190.74 0.39 ;
      LAYER M3 ;
      RECT 190.6 0.0 190.74 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[24]
  PIN DYA[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 387.19 0.0 387.33 0.39 ;
      LAYER M2 ;
      RECT 387.19 0.0 387.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[55]
  PIN DYA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 189.85 0.0 189.99 0.39 ;
      LAYER M1 ;
      RECT 189.85 0.0 189.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[24]
  PIN TDA[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 387.74 0.0 387.88 0.39 ;
      LAYER M4 ;
      RECT 387.74 0.0 387.88 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[55]
  PIN TDA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 189.3 0.0 189.44 0.39 ;
      LAYER M3 ;
      RECT 189.3 0.0 189.44 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[24]
  PIN TQA[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 387.98 0.0 388.12 0.39 ;
      LAYER M4 ;
      RECT 387.98 0.0 388.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[55]
  PIN TQA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 189.06 0.0 189.2 0.39 ;
      LAYER M3 ;
      RECT 189.06 0.0 189.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[24]
  PIN TQB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 388.55 0.0 388.69 0.39 ;
      LAYER M4 ;
      RECT 388.55 0.0 388.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[56]
  PIN TQB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 188.49 0.0 188.63 0.39 ;
      LAYER M3 ;
      RECT 188.49 0.0 188.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[23]
  PIN TDB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 388.79 0.0 388.93 0.39 ;
      LAYER M4 ;
      RECT 388.79 0.0 388.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[56]
  PIN TDB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 188.25 0.0 188.39 0.39 ;
      LAYER M3 ;
      RECT 188.25 0.0 188.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[23]
  PIN DYB[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 389.34 0.0 389.48 0.39 ;
      LAYER M2 ;
      RECT 389.34 0.0 389.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[56]
  PIN DYB[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 187.7 0.0 187.84 0.39 ;
      LAYER M1 ;
      RECT 187.7 0.0 187.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[23]
  PIN QB[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 390.09 0.0 390.23 0.39 ;
      LAYER M4 ;
      RECT 390.09 0.0 390.23 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[56]
  PIN QB[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 186.95 0.0 187.09 0.39 ;
      LAYER M3 ;
      RECT 186.95 0.0 187.09 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[23]
  PIN AYB[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 390.26 0.0 390.4 0.39 ;
      LAYER M2 ;
      RECT 390.26 0.0 390.4 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[9]
  PIN AYA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 186.78 0.0 186.92 0.39 ;
      LAYER M1 ;
      RECT 186.78 0.0 186.92 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[9]
  PIN DB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 391.08 0.0 391.22 0.39 ;
      LAYER M4 ;
      RECT 391.08 0.0 391.22 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[56]
  PIN DB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 185.96 0.0 186.1 0.39 ;
      LAYER M3 ;
      RECT 185.96 0.0 186.1 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[23]
  PIN AYB[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 391.115 0.0 391.255 0.39 ;
      LAYER M2 ;
      RECT 391.115 0.0 391.255 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYB[10]
  PIN AYA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 185.92 0.0 186.06 0.39 ;
      LAYER M1 ;
      RECT 185.92 0.0 186.06 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END AYA[10]
  PIN DA[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 391.65 0.0 391.79 0.39 ;
      LAYER M4 ;
      RECT 391.65 0.0 391.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[56]
  PIN DA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 185.39 0.0 185.53 0.39 ;
      LAYER M3 ;
      RECT 185.39 0.0 185.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[23]
  PIN QA[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 392.64 0.0 392.78 0.39 ;
      LAYER M4 ;
      RECT 392.64 0.0 392.78 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[56]
  PIN QA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 184.4 0.0 184.54 0.39 ;
      LAYER M3 ;
      RECT 184.4 0.0 184.54 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[23]
  PIN TAB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 392.75 0.0 392.89 0.39 ;
      LAYER M2 ;
      RECT 392.75 0.0 392.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[9]
  PIN TAA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 184.26 0.0 184.4 0.39 ;
      LAYER M1 ;
      RECT 184.26 0.0 184.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[9]
  PIN DYA[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 393.39 0.0 393.53 0.39 ;
      LAYER M2 ;
      RECT 393.39 0.0 393.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[56]
  PIN DYA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 183.65 0.0 183.79 0.39 ;
      LAYER M1 ;
      RECT 183.65 0.0 183.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[23]
  PIN TAB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 393.655 0.0 393.795 0.39 ;
      LAYER M2 ;
      RECT 393.655 0.0 393.795 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAB[10]
  PIN TAA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 183.365 0.0 183.505 0.39 ;
      LAYER M1 ;
      RECT 183.365 0.0 183.505 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TAA[10]
  PIN TDA[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 393.94 0.0 394.08 0.39 ;
      LAYER M4 ;
      RECT 393.94 0.0 394.08 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[56]
  PIN TDA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 183.1 0.0 183.24 0.39 ;
      LAYER M3 ;
      RECT 183.1 0.0 183.24 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[23]
  PIN TQA[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 394.18 0.0 394.32 0.39 ;
      LAYER M4 ;
      RECT 394.18 0.0 394.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[56]
  PIN TQA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 182.86 0.0 183.0 0.39 ;
      LAYER M3 ;
      RECT 182.86 0.0 183.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[23]
  PIN AB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 394.335 0.0 394.475 0.39 ;
      LAYER M2 ;
      RECT 394.335 0.0 394.475 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[10]
  PIN AA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 182.445 0.0 182.585 0.39 ;
      LAYER M1 ;
      RECT 182.445 0.0 182.585 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[10]
  PIN AB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 394.675 0.0 394.815 0.39 ;
      LAYER M2 ;
      RECT 394.675 0.0 394.815 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AB[9]
  PIN TQB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 182.29 0.0 182.43 0.39 ;
      LAYER M3 ;
      RECT 182.29 0.0 182.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[22]
  PIN TQB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 394.75 0.0 394.89 0.39 ;
      LAYER M4 ;
      RECT 394.75 0.0 394.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[57]
  PIN TDB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 182.05 0.0 182.19 0.39 ;
      LAYER M3 ;
      RECT 182.05 0.0 182.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[22]
  PIN TDB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 394.99 0.0 395.13 0.39 ;
      LAYER M4 ;
      RECT 394.99 0.0 395.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[57]
  PIN AA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 181.785 0.0 181.925 0.39 ;
      LAYER M1 ;
      RECT 181.785 0.0 181.925 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END AA[9]
  PIN CENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 395.24 0.0 395.38 0.39 ;
      LAYER M2 ;
      RECT 395.24 0.0 395.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END CENB
  PIN DYB[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 181.5 0.0 181.64 0.39 ;
      LAYER M1 ;
      RECT 181.5 0.0 181.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[22]
  PIN DYB[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 395.54 0.0 395.68 0.39 ;
      LAYER M2 ;
      RECT 395.54 0.0 395.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[57]
  PIN CENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 181.0 0.0 181.14 0.39 ;
      LAYER M1 ;
      RECT 181.0 0.0 181.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END CENA
  PIN WENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 396.24 0.0 396.38 0.39 ;
      LAYER M2 ;
      RECT 396.24 0.0 396.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END WENB
  PIN QB[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 180.75 0.0 180.89 0.39 ;
      LAYER M3 ;
      RECT 180.75 0.0 180.89 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[22]
  PIN QB[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 396.29 0.0 396.43 0.39 ;
      LAYER M4 ;
      RECT 396.29 0.0 396.43 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[57]
  PIN WENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 180.635 0.0 180.775 0.39 ;
      LAYER M1 ;
      RECT 180.635 0.0 180.775 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END WENA
  PIN TCENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 396.51 0.0 396.65 0.39 ;
      LAYER M2 ;
      RECT 396.51 0.0 396.65 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TCENB
  PIN DB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 179.76 0.0 179.9 0.39 ;
      LAYER M3 ;
      RECT 179.76 0.0 179.9 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[22]
  PIN DB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 397.28 0.0 397.42 0.39 ;
      LAYER M4 ;
      RECT 397.28 0.0 397.42 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[57]
  PIN TCENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 179.685 0.0 179.825 0.39 ;
      LAYER M1 ;
      RECT 179.685 0.0 179.825 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TCENA
  PIN TWENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 397.44 0.0 397.58 0.39 ;
      LAYER M2 ;
      RECT 397.44 0.0 397.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TWENB
  PIN TWENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 179.335 0.0 179.475 0.39 ;
      LAYER M1 ;
      RECT 179.335 0.0 179.475 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TWENA
  PIN DA[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 397.85 0.0 397.99 0.39 ;
      LAYER M4 ;
      RECT 397.85 0.0 397.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[57]
  PIN DA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 179.19 0.0 179.33 0.39 ;
      LAYER M3 ;
      RECT 179.19 0.0 179.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[22]
  PIN QA[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 398.84 0.0 398.98 0.39 ;
      LAYER M4 ;
      RECT 398.84 0.0 398.98 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[57]
  PIN QA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 178.2 0.0 178.34 0.39 ;
      LAYER M3 ;
      RECT 178.2 0.0 178.34 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[22]
  PIN DYA[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 399.59 0.0 399.73 0.39 ;
      LAYER M2 ;
      RECT 399.59 0.0 399.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[57]
  PIN DYA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 177.45 0.0 177.59 0.39 ;
      LAYER M1 ;
      RECT 177.45 0.0 177.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[22]
  PIN CENYB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 399.875 0.0 400.015 0.39 ;
      LAYER M2 ;
      RECT 399.875 0.0 400.015 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END CENYB
  PIN CENYA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 177.155 0.0 177.295 0.39 ;
      LAYER M1 ;
      RECT 177.155 0.0 177.295 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END CENYA
  PIN TDA[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 400.14 0.0 400.28 0.39 ;
      LAYER M4 ;
      RECT 400.14 0.0 400.28 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[57]
  PIN TDA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 176.9 0.0 177.04 0.39 ;
      LAYER M3 ;
      RECT 176.9 0.0 177.04 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[22]
  PIN TQA[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 400.38 0.0 400.52 0.39 ;
      LAYER M4 ;
      RECT 400.38 0.0 400.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[57]
  PIN TQA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 176.66 0.0 176.8 0.39 ;
      LAYER M3 ;
      RECT 176.66 0.0 176.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[22]
  PIN WENYB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 400.42 0.0 400.56 0.39 ;
      LAYER M2 ;
      RECT 400.42 0.0 400.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END WENYB
  PIN WENYA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 176.62 0.0 176.76 0.39 ;
      LAYER M1 ;
      RECT 176.62 0.0 176.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END WENYA
  PIN TQB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 400.98 0.0 401.12 0.39 ;
      LAYER M4 ;
      RECT 400.98 0.0 401.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[58]
  PIN TQB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 176.06 0.0 176.2 0.39 ;
      LAYER M3 ;
      RECT 176.06 0.0 176.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[21]
  PIN TDB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 401.23 0.0 401.37 0.39 ;
      LAYER M4 ;
      RECT 401.23 0.0 401.37 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[58]
  PIN TDB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 175.81 0.0 175.95 0.39 ;
      LAYER M3 ;
      RECT 175.81 0.0 175.95 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[21]
  PIN DYB[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 401.72 0.0 401.86 0.39 ;
      LAYER M2 ;
      RECT 401.72 0.0 401.86 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[58]
  PIN DYB[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 175.32 0.0 175.46 0.39 ;
      LAYER M1 ;
      RECT 175.32 0.0 175.46 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[21]
  PIN QB[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 402.49 0.0 402.63 0.39 ;
      LAYER M4 ;
      RECT 402.49 0.0 402.63 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[58]
  PIN QB[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 174.55 0.0 174.69 0.39 ;
      LAYER M3 ;
      RECT 174.55 0.0 174.69 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[21]
  PIN DB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 403.48 0.0 403.62 0.39 ;
      LAYER M4 ;
      RECT 403.48 0.0 403.62 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[58]
  PIN DB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 173.56 0.0 173.7 0.39 ;
      LAYER M3 ;
      RECT 173.56 0.0 173.7 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[21]
  PIN DA[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 404.05 0.0 404.19 0.39 ;
      LAYER M4 ;
      RECT 404.05 0.0 404.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[58]
  PIN DA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 172.99 0.0 173.13 0.39 ;
      LAYER M3 ;
      RECT 172.99 0.0 173.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[21]
  PIN QA[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 405.04 0.0 405.18 0.39 ;
      LAYER M4 ;
      RECT 405.04 0.0 405.18 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[58]
  PIN QA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 172.0 0.0 172.14 0.39 ;
      LAYER M3 ;
      RECT 172.0 0.0 172.14 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[21]
  PIN DYA[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 405.81 0.0 405.95 0.39 ;
      LAYER M2 ;
      RECT 405.81 0.0 405.95 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[58]
  PIN DYA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 171.23 0.0 171.37 0.39 ;
      LAYER M1 ;
      RECT 171.23 0.0 171.37 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[21]
  PIN TDA[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 406.305 0.0 406.445 0.39 ;
      LAYER M4 ;
      RECT 406.305 0.0 406.445 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[58]
  PIN TDA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 170.735 0.0 170.875 0.39 ;
      LAYER M3 ;
      RECT 170.735 0.0 170.875 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[21]
  PIN TQA[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 406.59 0.0 406.73 0.39 ;
      LAYER M4 ;
      RECT 406.59 0.0 406.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[58]
  PIN TQA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 170.45 0.0 170.59 0.39 ;
      LAYER M3 ;
      RECT 170.45 0.0 170.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[21]
  PIN TQB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 407.18 0.0 407.32 0.39 ;
      LAYER M4 ;
      RECT 407.18 0.0 407.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[59]
  PIN TQB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 169.86 0.0 170.0 0.39 ;
      LAYER M3 ;
      RECT 169.86 0.0 170.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[20]
  PIN TDB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 407.43 0.0 407.57 0.39 ;
      LAYER M4 ;
      RECT 407.43 0.0 407.57 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[59]
  PIN TDB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 169.61 0.0 169.75 0.39 ;
      LAYER M3 ;
      RECT 169.61 0.0 169.75 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[20]
  PIN DYB[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 407.92 0.0 408.06 0.39 ;
      LAYER M2 ;
      RECT 407.92 0.0 408.06 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[59]
  PIN DYB[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 169.12 0.0 169.26 0.39 ;
      LAYER M1 ;
      RECT 169.12 0.0 169.26 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[20]
  PIN QB[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 408.69 0.0 408.83 0.39 ;
      LAYER M4 ;
      RECT 408.69 0.0 408.83 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[59]
  PIN QB[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 168.35 0.0 168.49 0.39 ;
      LAYER M3 ;
      RECT 168.35 0.0 168.49 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[20]
  PIN DB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 409.68 0.0 409.82 0.39 ;
      LAYER M4 ;
      RECT 409.68 0.0 409.82 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[59]
  PIN DB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 167.36 0.0 167.5 0.39 ;
      LAYER M3 ;
      RECT 167.36 0.0 167.5 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[20]
  PIN DA[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 410.25 0.0 410.39 0.39 ;
      LAYER M4 ;
      RECT 410.25 0.0 410.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[59]
  PIN DA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 166.79 0.0 166.93 0.39 ;
      LAYER M3 ;
      RECT 166.79 0.0 166.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[20]
  PIN QA[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 411.24 0.0 411.38 0.39 ;
      LAYER M4 ;
      RECT 411.24 0.0 411.38 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[59]
  PIN QA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 165.8 0.0 165.94 0.39 ;
      LAYER M3 ;
      RECT 165.8 0.0 165.94 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[20]
  PIN DYA[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 412.01 0.0 412.15 0.39 ;
      LAYER M2 ;
      RECT 412.01 0.0 412.15 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[59]
  PIN DYA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 165.03 0.0 165.17 0.39 ;
      LAYER M1 ;
      RECT 165.03 0.0 165.17 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[20]
  PIN TDA[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 412.505 0.0 412.645 0.39 ;
      LAYER M4 ;
      RECT 412.505 0.0 412.645 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[59]
  PIN TDA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 164.535 0.0 164.675 0.39 ;
      LAYER M3 ;
      RECT 164.535 0.0 164.675 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[20]
  PIN TQA[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 412.79 0.0 412.93 0.39 ;
      LAYER M4 ;
      RECT 412.79 0.0 412.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[59]
  PIN TQA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 164.25 0.0 164.39 0.39 ;
      LAYER M3 ;
      RECT 164.25 0.0 164.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[20]
  PIN TQB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 452.59 0.0 452.73 0.39 ;
      LAYER M4 ;
      RECT 452.59 0.0 452.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[60]
  PIN TQB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 124.45 0.0 124.59 0.39 ;
      LAYER M3 ;
      RECT 124.45 0.0 124.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[19]
  PIN TDB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 452.84 0.0 452.98 0.39 ;
      LAYER M4 ;
      RECT 452.84 0.0 452.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[60]
  PIN TDB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 124.2 0.0 124.34 0.39 ;
      LAYER M3 ;
      RECT 124.2 0.0 124.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[19]
  PIN DYB[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 453.33 0.0 453.47 0.39 ;
      LAYER M2 ;
      RECT 453.33 0.0 453.47 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[60]
  PIN DYB[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 123.71 0.0 123.85 0.39 ;
      LAYER M1 ;
      RECT 123.71 0.0 123.85 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[19]
  PIN QB[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 454.1 0.0 454.24 0.39 ;
      LAYER M4 ;
      RECT 454.1 0.0 454.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[60]
  PIN QB[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 122.94 0.0 123.08 0.39 ;
      LAYER M3 ;
      RECT 122.94 0.0 123.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[19]
  PIN DB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 455.09 0.0 455.23 0.39 ;
      LAYER M4 ;
      RECT 455.09 0.0 455.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[60]
  PIN DB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 121.95 0.0 122.09 0.39 ;
      LAYER M3 ;
      RECT 121.95 0.0 122.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[19]
  PIN DA[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 455.66 0.0 455.8 0.39 ;
      LAYER M4 ;
      RECT 455.66 0.0 455.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[60]
  PIN DA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 121.38 0.0 121.52 0.39 ;
      LAYER M3 ;
      RECT 121.38 0.0 121.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[19]
  PIN QA[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 456.65 0.0 456.79 0.39 ;
      LAYER M4 ;
      RECT 456.65 0.0 456.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[60]
  PIN QA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 120.39 0.0 120.53 0.39 ;
      LAYER M3 ;
      RECT 120.39 0.0 120.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[19]
  PIN DYA[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 457.42 0.0 457.56 0.39 ;
      LAYER M2 ;
      RECT 457.42 0.0 457.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[60]
  PIN DYA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 119.62 0.0 119.76 0.39 ;
      LAYER M1 ;
      RECT 119.62 0.0 119.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[19]
  PIN TDA[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 457.915 0.0 458.055 0.39 ;
      LAYER M4 ;
      RECT 457.915 0.0 458.055 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[60]
  PIN TDA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 119.125 0.0 119.265 0.39 ;
      LAYER M3 ;
      RECT 119.125 0.0 119.265 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[19]
  PIN TQA[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 458.2 0.0 458.34 0.39 ;
      LAYER M4 ;
      RECT 458.2 0.0 458.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[60]
  PIN TQA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 118.84 0.0 118.98 0.39 ;
      LAYER M3 ;
      RECT 118.84 0.0 118.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[19]
  PIN TQB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 458.79 0.0 458.93 0.39 ;
      LAYER M4 ;
      RECT 458.79 0.0 458.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[61]
  PIN TQB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 118.25 0.0 118.39 0.39 ;
      LAYER M3 ;
      RECT 118.25 0.0 118.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[18]
  PIN TDB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 459.04 0.0 459.18 0.39 ;
      LAYER M4 ;
      RECT 459.04 0.0 459.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[61]
  PIN TDB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 118.0 0.0 118.14 0.39 ;
      LAYER M3 ;
      RECT 118.0 0.0 118.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[18]
  PIN DYB[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 459.53 0.0 459.67 0.39 ;
      LAYER M2 ;
      RECT 459.53 0.0 459.67 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[61]
  PIN DYB[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 117.51 0.0 117.65 0.39 ;
      LAYER M1 ;
      RECT 117.51 0.0 117.65 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[18]
  PIN QB[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 460.3 0.0 460.44 0.39 ;
      LAYER M4 ;
      RECT 460.3 0.0 460.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[61]
  PIN QB[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 116.74 0.0 116.88 0.39 ;
      LAYER M3 ;
      RECT 116.74 0.0 116.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[18]
  PIN DB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 461.29 0.0 461.43 0.39 ;
      LAYER M4 ;
      RECT 461.29 0.0 461.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[61]
  PIN DB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 115.75 0.0 115.89 0.39 ;
      LAYER M3 ;
      RECT 115.75 0.0 115.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[18]
  PIN DA[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 461.86 0.0 462.0 0.39 ;
      LAYER M4 ;
      RECT 461.86 0.0 462.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[61]
  PIN DA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 115.18 0.0 115.32 0.39 ;
      LAYER M3 ;
      RECT 115.18 0.0 115.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[18]
  PIN QA[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 462.85 0.0 462.99 0.39 ;
      LAYER M4 ;
      RECT 462.85 0.0 462.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[61]
  PIN QA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 114.19 0.0 114.33 0.39 ;
      LAYER M3 ;
      RECT 114.19 0.0 114.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[18]
  PIN DYA[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 463.62 0.0 463.76 0.39 ;
      LAYER M2 ;
      RECT 463.62 0.0 463.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[61]
  PIN DYA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 113.42 0.0 113.56 0.39 ;
      LAYER M1 ;
      RECT 113.42 0.0 113.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[18]
  PIN TDA[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 464.115 0.0 464.255 0.39 ;
      LAYER M4 ;
      RECT 464.115 0.0 464.255 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[61]
  PIN TDA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 112.925 0.0 113.065 0.39 ;
      LAYER M3 ;
      RECT 112.925 0.0 113.065 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[18]
  PIN TQA[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 464.4 0.0 464.54 0.39 ;
      LAYER M4 ;
      RECT 464.4 0.0 464.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[61]
  PIN TQA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 112.64 0.0 112.78 0.39 ;
      LAYER M3 ;
      RECT 112.64 0.0 112.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[18]
  PIN TQB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 464.99 0.0 465.13 0.39 ;
      LAYER M4 ;
      RECT 464.99 0.0 465.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[62]
  PIN TQB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 112.05 0.0 112.19 0.39 ;
      LAYER M3 ;
      RECT 112.05 0.0 112.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[17]
  PIN TDB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 465.24 0.0 465.38 0.39 ;
      LAYER M4 ;
      RECT 465.24 0.0 465.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[62]
  PIN TDB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 111.8 0.0 111.94 0.39 ;
      LAYER M3 ;
      RECT 111.8 0.0 111.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[17]
  PIN DYB[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 465.73 0.0 465.87 0.39 ;
      LAYER M2 ;
      RECT 465.73 0.0 465.87 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[62]
  PIN DYB[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 111.31 0.0 111.45 0.39 ;
      LAYER M1 ;
      RECT 111.31 0.0 111.45 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[17]
  PIN QB[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 466.5 0.0 466.64 0.39 ;
      LAYER M4 ;
      RECT 466.5 0.0 466.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[62]
  PIN QB[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 110.54 0.0 110.68 0.39 ;
      LAYER M3 ;
      RECT 110.54 0.0 110.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[17]
  PIN DB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 467.49 0.0 467.63 0.39 ;
      LAYER M4 ;
      RECT 467.49 0.0 467.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[62]
  PIN DB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 109.55 0.0 109.69 0.39 ;
      LAYER M3 ;
      RECT 109.55 0.0 109.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[17]
  PIN DA[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 468.06 0.0 468.2 0.39 ;
      LAYER M4 ;
      RECT 468.06 0.0 468.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[62]
  PIN DA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 108.98 0.0 109.12 0.39 ;
      LAYER M3 ;
      RECT 108.98 0.0 109.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[17]
  PIN QA[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 469.05 0.0 469.19 0.39 ;
      LAYER M4 ;
      RECT 469.05 0.0 469.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[62]
  PIN QA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 107.99 0.0 108.13 0.39 ;
      LAYER M3 ;
      RECT 107.99 0.0 108.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[17]
  PIN DYA[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 469.82 0.0 469.96 0.39 ;
      LAYER M2 ;
      RECT 469.82 0.0 469.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[62]
  PIN DYA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 107.22 0.0 107.36 0.39 ;
      LAYER M1 ;
      RECT 107.22 0.0 107.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[17]
  PIN TDA[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 470.315 0.0 470.455 0.39 ;
      LAYER M4 ;
      RECT 470.315 0.0 470.455 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[62]
  PIN TDA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 106.725 0.0 106.865 0.39 ;
      LAYER M3 ;
      RECT 106.725 0.0 106.865 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[17]
  PIN TQA[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 470.6 0.0 470.74 0.39 ;
      LAYER M4 ;
      RECT 470.6 0.0 470.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[62]
  PIN TQA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 106.44 0.0 106.58 0.39 ;
      LAYER M3 ;
      RECT 106.44 0.0 106.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[17]
  PIN TQB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 471.19 0.0 471.33 0.39 ;
      LAYER M4 ;
      RECT 471.19 0.0 471.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[63]
  PIN TQB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 105.85 0.0 105.99 0.39 ;
      LAYER M3 ;
      RECT 105.85 0.0 105.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[16]
  PIN TDB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 471.44 0.0 471.58 0.39 ;
      LAYER M4 ;
      RECT 471.44 0.0 471.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[63]
  PIN TDB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 105.6 0.0 105.74 0.39 ;
      LAYER M3 ;
      RECT 105.6 0.0 105.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[16]
  PIN DYB[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 471.93 0.0 472.07 0.39 ;
      LAYER M2 ;
      RECT 471.93 0.0 472.07 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[63]
  PIN DYB[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 105.11 0.0 105.25 0.39 ;
      LAYER M1 ;
      RECT 105.11 0.0 105.25 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[16]
  PIN QB[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 472.7 0.0 472.84 0.39 ;
      LAYER M4 ;
      RECT 472.7 0.0 472.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[63]
  PIN QB[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 104.34 0.0 104.48 0.39 ;
      LAYER M3 ;
      RECT 104.34 0.0 104.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[16]
  PIN DB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 473.69 0.0 473.83 0.39 ;
      LAYER M4 ;
      RECT 473.69 0.0 473.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[63]
  PIN DB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 103.35 0.0 103.49 0.39 ;
      LAYER M3 ;
      RECT 103.35 0.0 103.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[16]
  PIN DA[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 474.26 0.0 474.4 0.39 ;
      LAYER M4 ;
      RECT 474.26 0.0 474.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[63]
  PIN DA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 102.78 0.0 102.92 0.39 ;
      LAYER M3 ;
      RECT 102.78 0.0 102.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[16]
  PIN QA[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 475.25 0.0 475.39 0.39 ;
      LAYER M4 ;
      RECT 475.25 0.0 475.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[63]
  PIN QA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 101.79 0.0 101.93 0.39 ;
      LAYER M3 ;
      RECT 101.79 0.0 101.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[16]
  PIN DYA[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 476.02 0.0 476.16 0.39 ;
      LAYER M2 ;
      RECT 476.02 0.0 476.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[63]
  PIN DYA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 101.02 0.0 101.16 0.39 ;
      LAYER M1 ;
      RECT 101.02 0.0 101.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[16]
  PIN TDA[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 476.515 0.0 476.655 0.39 ;
      LAYER M4 ;
      RECT 476.515 0.0 476.655 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[63]
  PIN TDA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 100.525 0.0 100.665 0.39 ;
      LAYER M3 ;
      RECT 100.525 0.0 100.665 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[16]
  PIN TQA[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 476.8 0.0 476.94 0.39 ;
      LAYER M4 ;
      RECT 476.8 0.0 476.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[63]
  PIN TQA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 100.24 0.0 100.38 0.39 ;
      LAYER M3 ;
      RECT 100.24 0.0 100.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[16]
  PIN TQB[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 477.39 0.0 477.53 0.39 ;
      LAYER M4 ;
      RECT 477.39 0.0 477.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[64]
  PIN TQB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 99.65 0.0 99.79 0.39 ;
      LAYER M3 ;
      RECT 99.65 0.0 99.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[15]
  PIN TDB[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 477.64 0.0 477.78 0.39 ;
      LAYER M4 ;
      RECT 477.64 0.0 477.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[64]
  PIN TDB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 99.4 0.0 99.54 0.39 ;
      LAYER M3 ;
      RECT 99.4 0.0 99.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[15]
  PIN DYB[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 478.13 0.0 478.27 0.39 ;
      LAYER M2 ;
      RECT 478.13 0.0 478.27 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[64]
  PIN DYB[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 98.91 0.0 99.05 0.39 ;
      LAYER M1 ;
      RECT 98.91 0.0 99.05 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[15]
  PIN QB[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 478.9 0.0 479.04 0.39 ;
      LAYER M4 ;
      RECT 478.9 0.0 479.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[64]
  PIN QB[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 98.14 0.0 98.28 0.39 ;
      LAYER M3 ;
      RECT 98.14 0.0 98.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[15]
  PIN DB[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 479.89 0.0 480.03 0.39 ;
      LAYER M4 ;
      RECT 479.89 0.0 480.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[64]
  PIN DB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 97.15 0.0 97.29 0.39 ;
      LAYER M3 ;
      RECT 97.15 0.0 97.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[15]
  PIN DA[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 480.46 0.0 480.6 0.39 ;
      LAYER M4 ;
      RECT 480.46 0.0 480.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[64]
  PIN DA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 96.58 0.0 96.72 0.39 ;
      LAYER M3 ;
      RECT 96.58 0.0 96.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[15]
  PIN QA[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 481.45 0.0 481.59 0.39 ;
      LAYER M4 ;
      RECT 481.45 0.0 481.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[64]
  PIN QA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 95.59 0.0 95.73 0.39 ;
      LAYER M3 ;
      RECT 95.59 0.0 95.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[15]
  PIN DYA[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 482.22 0.0 482.36 0.39 ;
      LAYER M2 ;
      RECT 482.22 0.0 482.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[64]
  PIN DYA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 94.82 0.0 94.96 0.39 ;
      LAYER M1 ;
      RECT 94.82 0.0 94.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[15]
  PIN TDA[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 482.715 0.0 482.855 0.39 ;
      LAYER M4 ;
      RECT 482.715 0.0 482.855 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[64]
  PIN TDA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 94.325 0.0 94.465 0.39 ;
      LAYER M3 ;
      RECT 94.325 0.0 94.465 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[15]
  PIN TQA[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 483.0 0.0 483.14 0.39 ;
      LAYER M4 ;
      RECT 483.0 0.0 483.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[64]
  PIN TQA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 94.04 0.0 94.18 0.39 ;
      LAYER M3 ;
      RECT 94.04 0.0 94.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[15]
  PIN TQB[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 483.59 0.0 483.73 0.39 ;
      LAYER M4 ;
      RECT 483.59 0.0 483.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[65]
  PIN TQB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 93.45 0.0 93.59 0.39 ;
      LAYER M3 ;
      RECT 93.45 0.0 93.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[14]
  PIN TDB[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 483.84 0.0 483.98 0.39 ;
      LAYER M4 ;
      RECT 483.84 0.0 483.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[65]
  PIN TDB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 93.2 0.0 93.34 0.39 ;
      LAYER M3 ;
      RECT 93.2 0.0 93.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[14]
  PIN DYB[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 484.33 0.0 484.47 0.39 ;
      LAYER M2 ;
      RECT 484.33 0.0 484.47 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[65]
  PIN DYB[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 92.71 0.0 92.85 0.39 ;
      LAYER M1 ;
      RECT 92.71 0.0 92.85 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[14]
  PIN QB[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 485.1 0.0 485.24 0.39 ;
      LAYER M4 ;
      RECT 485.1 0.0 485.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[65]
  PIN QB[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 91.94 0.0 92.08 0.39 ;
      LAYER M3 ;
      RECT 91.94 0.0 92.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[14]
  PIN DB[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 486.09 0.0 486.23 0.39 ;
      LAYER M4 ;
      RECT 486.09 0.0 486.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[65]
  PIN DB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 90.95 0.0 91.09 0.39 ;
      LAYER M3 ;
      RECT 90.95 0.0 91.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[14]
  PIN DA[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 486.66 0.0 486.8 0.39 ;
      LAYER M4 ;
      RECT 486.66 0.0 486.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[65]
  PIN DA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 90.38 0.0 90.52 0.39 ;
      LAYER M3 ;
      RECT 90.38 0.0 90.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[14]
  PIN QA[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 487.65 0.0 487.79 0.39 ;
      LAYER M4 ;
      RECT 487.65 0.0 487.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[65]
  PIN QA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 89.39 0.0 89.53 0.39 ;
      LAYER M3 ;
      RECT 89.39 0.0 89.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[14]
  PIN DYA[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 488.42 0.0 488.56 0.39 ;
      LAYER M2 ;
      RECT 488.42 0.0 488.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[65]
  PIN DYA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 88.62 0.0 88.76 0.39 ;
      LAYER M1 ;
      RECT 88.62 0.0 88.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[14]
  PIN TDA[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 488.915 0.0 489.055 0.39 ;
      LAYER M4 ;
      RECT 488.915 0.0 489.055 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[65]
  PIN TDA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 88.125 0.0 88.265 0.39 ;
      LAYER M3 ;
      RECT 88.125 0.0 88.265 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[14]
  PIN TQA[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 489.2 0.0 489.34 0.39 ;
      LAYER M4 ;
      RECT 489.2 0.0 489.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[65]
  PIN TQA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 87.84 0.0 87.98 0.39 ;
      LAYER M3 ;
      RECT 87.84 0.0 87.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[14]
  PIN TQB[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 489.79 0.0 489.93 0.39 ;
      LAYER M4 ;
      RECT 489.79 0.0 489.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[66]
  PIN TQB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 87.25 0.0 87.39 0.39 ;
      LAYER M3 ;
      RECT 87.25 0.0 87.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[13]
  PIN TDB[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 490.04 0.0 490.18 0.39 ;
      LAYER M4 ;
      RECT 490.04 0.0 490.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[66]
  PIN TDB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 87.0 0.0 87.14 0.39 ;
      LAYER M3 ;
      RECT 87.0 0.0 87.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[13]
  PIN DYB[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 490.53 0.0 490.67 0.39 ;
      LAYER M2 ;
      RECT 490.53 0.0 490.67 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[66]
  PIN DYB[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 86.51 0.0 86.65 0.39 ;
      LAYER M1 ;
      RECT 86.51 0.0 86.65 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[13]
  PIN QB[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 491.3 0.0 491.44 0.39 ;
      LAYER M4 ;
      RECT 491.3 0.0 491.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[66]
  PIN QB[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 85.74 0.0 85.88 0.39 ;
      LAYER M3 ;
      RECT 85.74 0.0 85.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[13]
  PIN DB[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 492.29 0.0 492.43 0.39 ;
      LAYER M4 ;
      RECT 492.29 0.0 492.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[66]
  PIN DB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 84.75 0.0 84.89 0.39 ;
      LAYER M3 ;
      RECT 84.75 0.0 84.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[13]
  PIN DA[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 492.86 0.0 493.0 0.39 ;
      LAYER M4 ;
      RECT 492.86 0.0 493.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[66]
  PIN DA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 84.18 0.0 84.32 0.39 ;
      LAYER M3 ;
      RECT 84.18 0.0 84.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[13]
  PIN QA[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 493.85 0.0 493.99 0.39 ;
      LAYER M4 ;
      RECT 493.85 0.0 493.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[66]
  PIN QA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 83.19 0.0 83.33 0.39 ;
      LAYER M3 ;
      RECT 83.19 0.0 83.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[13]
  PIN DYA[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 494.62 0.0 494.76 0.39 ;
      LAYER M2 ;
      RECT 494.62 0.0 494.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[66]
  PIN DYA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 82.42 0.0 82.56 0.39 ;
      LAYER M1 ;
      RECT 82.42 0.0 82.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[13]
  PIN TDA[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 495.115 0.0 495.255 0.39 ;
      LAYER M4 ;
      RECT 495.115 0.0 495.255 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[66]
  PIN TDA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 81.925 0.0 82.065 0.39 ;
      LAYER M3 ;
      RECT 81.925 0.0 82.065 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[13]
  PIN TQA[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 495.4 0.0 495.54 0.39 ;
      LAYER M4 ;
      RECT 495.4 0.0 495.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[66]
  PIN TQA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 81.64 0.0 81.78 0.39 ;
      LAYER M3 ;
      RECT 81.64 0.0 81.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[13]
  PIN TQB[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 495.99 0.0 496.13 0.39 ;
      LAYER M4 ;
      RECT 495.99 0.0 496.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[67]
  PIN TQB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 81.05 0.0 81.19 0.39 ;
      LAYER M3 ;
      RECT 81.05 0.0 81.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[12]
  PIN TDB[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 496.24 0.0 496.38 0.39 ;
      LAYER M4 ;
      RECT 496.24 0.0 496.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[67]
  PIN TDB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 80.8 0.0 80.94 0.39 ;
      LAYER M3 ;
      RECT 80.8 0.0 80.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[12]
  PIN DYB[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 496.73 0.0 496.87 0.39 ;
      LAYER M2 ;
      RECT 496.73 0.0 496.87 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[67]
  PIN DYB[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 80.31 0.0 80.45 0.39 ;
      LAYER M1 ;
      RECT 80.31 0.0 80.45 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[12]
  PIN QB[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 497.5 0.0 497.64 0.39 ;
      LAYER M4 ;
      RECT 497.5 0.0 497.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[67]
  PIN QB[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 79.54 0.0 79.68 0.39 ;
      LAYER M3 ;
      RECT 79.54 0.0 79.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[12]
  PIN DB[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 498.49 0.0 498.63 0.39 ;
      LAYER M4 ;
      RECT 498.49 0.0 498.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[67]
  PIN DB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 78.55 0.0 78.69 0.39 ;
      LAYER M3 ;
      RECT 78.55 0.0 78.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[12]
  PIN DA[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 499.06 0.0 499.2 0.39 ;
      LAYER M4 ;
      RECT 499.06 0.0 499.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[67]
  PIN DA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 77.98 0.0 78.12 0.39 ;
      LAYER M3 ;
      RECT 77.98 0.0 78.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[12]
  PIN QA[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 500.05 0.0 500.19 0.39 ;
      LAYER M4 ;
      RECT 500.05 0.0 500.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[67]
  PIN QA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 76.99 0.0 77.13 0.39 ;
      LAYER M3 ;
      RECT 76.99 0.0 77.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[12]
  PIN DYA[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 500.82 0.0 500.96 0.39 ;
      LAYER M2 ;
      RECT 500.82 0.0 500.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[67]
  PIN DYA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 76.22 0.0 76.36 0.39 ;
      LAYER M1 ;
      RECT 76.22 0.0 76.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[12]
  PIN TDA[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 501.315 0.0 501.455 0.39 ;
      LAYER M4 ;
      RECT 501.315 0.0 501.455 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[67]
  PIN TDA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 75.725 0.0 75.865 0.39 ;
      LAYER M3 ;
      RECT 75.725 0.0 75.865 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[12]
  PIN TQA[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 501.6 0.0 501.74 0.39 ;
      LAYER M4 ;
      RECT 501.6 0.0 501.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[67]
  PIN TQA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 75.44 0.0 75.58 0.39 ;
      LAYER M3 ;
      RECT 75.44 0.0 75.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[12]
  PIN TQB[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 502.19 0.0 502.33 0.39 ;
      LAYER M4 ;
      RECT 502.19 0.0 502.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[68]
  PIN TQB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 74.85 0.0 74.99 0.39 ;
      LAYER M3 ;
      RECT 74.85 0.0 74.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[11]
  PIN TDB[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 502.44 0.0 502.58 0.39 ;
      LAYER M4 ;
      RECT 502.44 0.0 502.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[68]
  PIN TDB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 74.6 0.0 74.74 0.39 ;
      LAYER M3 ;
      RECT 74.6 0.0 74.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[11]
  PIN DYB[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 502.93 0.0 503.07 0.39 ;
      LAYER M2 ;
      RECT 502.93 0.0 503.07 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[68]
  PIN DYB[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 74.11 0.0 74.25 0.39 ;
      LAYER M1 ;
      RECT 74.11 0.0 74.25 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[11]
  PIN QB[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 503.7 0.0 503.84 0.39 ;
      LAYER M4 ;
      RECT 503.7 0.0 503.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[68]
  PIN QB[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 73.34 0.0 73.48 0.39 ;
      LAYER M3 ;
      RECT 73.34 0.0 73.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[11]
  PIN DB[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 504.69 0.0 504.83 0.39 ;
      LAYER M4 ;
      RECT 504.69 0.0 504.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[68]
  PIN DB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 72.35 0.0 72.49 0.39 ;
      LAYER M3 ;
      RECT 72.35 0.0 72.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[11]
  PIN DA[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 505.26 0.0 505.4 0.39 ;
      LAYER M4 ;
      RECT 505.26 0.0 505.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[68]
  PIN DA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 71.78 0.0 71.92 0.39 ;
      LAYER M3 ;
      RECT 71.78 0.0 71.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[11]
  PIN QA[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 506.25 0.0 506.39 0.39 ;
      LAYER M4 ;
      RECT 506.25 0.0 506.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[68]
  PIN QA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 70.79 0.0 70.93 0.39 ;
      LAYER M3 ;
      RECT 70.79 0.0 70.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[11]
  PIN DYA[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 507.02 0.0 507.16 0.39 ;
      LAYER M2 ;
      RECT 507.02 0.0 507.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[68]
  PIN DYA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 70.02 0.0 70.16 0.39 ;
      LAYER M1 ;
      RECT 70.02 0.0 70.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[11]
  PIN TDA[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 507.515 0.0 507.655 0.39 ;
      LAYER M4 ;
      RECT 507.515 0.0 507.655 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[68]
  PIN TDA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 69.525 0.0 69.665 0.39 ;
      LAYER M3 ;
      RECT 69.525 0.0 69.665 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[11]
  PIN TQA[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 507.8 0.0 507.94 0.39 ;
      LAYER M4 ;
      RECT 507.8 0.0 507.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[68]
  PIN TQA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 69.24 0.0 69.38 0.39 ;
      LAYER M3 ;
      RECT 69.24 0.0 69.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[11]
  PIN TQB[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 508.39 0.0 508.53 0.39 ;
      LAYER M4 ;
      RECT 508.39 0.0 508.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[69]
  PIN TQB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 68.65 0.0 68.79 0.39 ;
      LAYER M3 ;
      RECT 68.65 0.0 68.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[10]
  PIN TDB[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 508.64 0.0 508.78 0.39 ;
      LAYER M4 ;
      RECT 508.64 0.0 508.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[69]
  PIN TDB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 68.4 0.0 68.54 0.39 ;
      LAYER M3 ;
      RECT 68.4 0.0 68.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[10]
  PIN DYB[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 509.13 0.0 509.27 0.39 ;
      LAYER M2 ;
      RECT 509.13 0.0 509.27 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[69]
  PIN DYB[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 67.91 0.0 68.05 0.39 ;
      LAYER M1 ;
      RECT 67.91 0.0 68.05 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[10]
  PIN QB[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 509.9 0.0 510.04 0.39 ;
      LAYER M4 ;
      RECT 509.9 0.0 510.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[69]
  PIN QB[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 67.14 0.0 67.28 0.39 ;
      LAYER M3 ;
      RECT 67.14 0.0 67.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[10]
  PIN DB[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 510.89 0.0 511.03 0.39 ;
      LAYER M4 ;
      RECT 510.89 0.0 511.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[69]
  PIN DB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 66.15 0.0 66.29 0.39 ;
      LAYER M3 ;
      RECT 66.15 0.0 66.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[10]
  PIN DA[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 511.46 0.0 511.6 0.39 ;
      LAYER M4 ;
      RECT 511.46 0.0 511.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[69]
  PIN DA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 65.58 0.0 65.72 0.39 ;
      LAYER M3 ;
      RECT 65.58 0.0 65.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[10]
  PIN QA[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 512.45 0.0 512.59 0.39 ;
      LAYER M4 ;
      RECT 512.45 0.0 512.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[69]
  PIN QA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 64.59 0.0 64.73 0.39 ;
      LAYER M3 ;
      RECT 64.59 0.0 64.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[10]
  PIN DYA[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 513.22 0.0 513.36 0.39 ;
      LAYER M2 ;
      RECT 513.22 0.0 513.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[69]
  PIN DYA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 63.82 0.0 63.96 0.39 ;
      LAYER M1 ;
      RECT 63.82 0.0 63.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[10]
  PIN TDA[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 513.715 0.0 513.855 0.39 ;
      LAYER M4 ;
      RECT 513.715 0.0 513.855 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[69]
  PIN TDA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 63.325 0.0 63.465 0.39 ;
      LAYER M3 ;
      RECT 63.325 0.0 63.465 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[10]
  PIN TQA[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 514.0 0.0 514.14 0.39 ;
      LAYER M4 ;
      RECT 514.0 0.0 514.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[69]
  PIN TQA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 63.04 0.0 63.18 0.39 ;
      LAYER M3 ;
      RECT 63.04 0.0 63.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[10]
  PIN TQB[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 514.59 0.0 514.73 0.39 ;
      LAYER M4 ;
      RECT 514.59 0.0 514.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[70]
  PIN TQB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 62.45 0.0 62.59 0.39 ;
      LAYER M3 ;
      RECT 62.45 0.0 62.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[9]
  PIN TDB[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 514.84 0.0 514.98 0.39 ;
      LAYER M4 ;
      RECT 514.84 0.0 514.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[70]
  PIN TDB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 62.2 0.0 62.34 0.39 ;
      LAYER M3 ;
      RECT 62.2 0.0 62.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[9]
  PIN DYB[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 515.33 0.0 515.47 0.39 ;
      LAYER M2 ;
      RECT 515.33 0.0 515.47 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[70]
  PIN DYB[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 61.71 0.0 61.85 0.39 ;
      LAYER M1 ;
      RECT 61.71 0.0 61.85 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[9]
  PIN QB[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 516.1 0.0 516.24 0.39 ;
      LAYER M4 ;
      RECT 516.1 0.0 516.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[70]
  PIN QB[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 60.94 0.0 61.08 0.39 ;
      LAYER M3 ;
      RECT 60.94 0.0 61.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[9]
  PIN DB[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 517.09 0.0 517.23 0.39 ;
      LAYER M4 ;
      RECT 517.09 0.0 517.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[70]
  PIN DB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 59.95 0.0 60.09 0.39 ;
      LAYER M3 ;
      RECT 59.95 0.0 60.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[9]
  PIN DA[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 517.66 0.0 517.8 0.39 ;
      LAYER M4 ;
      RECT 517.66 0.0 517.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[70]
  PIN DA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 59.38 0.0 59.52 0.39 ;
      LAYER M3 ;
      RECT 59.38 0.0 59.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[9]
  PIN QA[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 518.65 0.0 518.79 0.39 ;
      LAYER M4 ;
      RECT 518.65 0.0 518.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[70]
  PIN QA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 58.39 0.0 58.53 0.39 ;
      LAYER M3 ;
      RECT 58.39 0.0 58.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[9]
  PIN DYA[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 519.42 0.0 519.56 0.39 ;
      LAYER M2 ;
      RECT 519.42 0.0 519.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[70]
  PIN DYA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 57.62 0.0 57.76 0.39 ;
      LAYER M1 ;
      RECT 57.62 0.0 57.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[9]
  PIN TDA[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 519.915 0.0 520.055 0.39 ;
      LAYER M4 ;
      RECT 519.915 0.0 520.055 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[70]
  PIN TDA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 57.125 0.0 57.265 0.39 ;
      LAYER M3 ;
      RECT 57.125 0.0 57.265 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[9]
  PIN TQA[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 520.2 0.0 520.34 0.39 ;
      LAYER M4 ;
      RECT 520.2 0.0 520.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[70]
  PIN TQA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 56.84 0.0 56.98 0.39 ;
      LAYER M3 ;
      RECT 56.84 0.0 56.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[9]
  PIN TQB[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 520.79 0.0 520.93 0.39 ;
      LAYER M4 ;
      RECT 520.79 0.0 520.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[71]
  PIN TQB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 56.25 0.0 56.39 0.39 ;
      LAYER M3 ;
      RECT 56.25 0.0 56.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[8]
  PIN TDB[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 521.04 0.0 521.18 0.39 ;
      LAYER M4 ;
      RECT 521.04 0.0 521.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[71]
  PIN TDB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 56.0 0.0 56.14 0.39 ;
      LAYER M3 ;
      RECT 56.0 0.0 56.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[8]
  PIN DYB[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 521.53 0.0 521.67 0.39 ;
      LAYER M2 ;
      RECT 521.53 0.0 521.67 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[71]
  PIN DYB[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 55.51 0.0 55.65 0.39 ;
      LAYER M1 ;
      RECT 55.51 0.0 55.65 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[8]
  PIN QB[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 522.3 0.0 522.44 0.39 ;
      LAYER M4 ;
      RECT 522.3 0.0 522.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[71]
  PIN QB[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 54.74 0.0 54.88 0.39 ;
      LAYER M3 ;
      RECT 54.74 0.0 54.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[8]
  PIN DB[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 523.29 0.0 523.43 0.39 ;
      LAYER M4 ;
      RECT 523.29 0.0 523.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[71]
  PIN DB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 53.75 0.0 53.89 0.39 ;
      LAYER M3 ;
      RECT 53.75 0.0 53.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[8]
  PIN DA[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 523.86 0.0 524.0 0.39 ;
      LAYER M4 ;
      RECT 523.86 0.0 524.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[71]
  PIN DA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 53.18 0.0 53.32 0.39 ;
      LAYER M3 ;
      RECT 53.18 0.0 53.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[8]
  PIN QA[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 524.85 0.0 524.99 0.39 ;
      LAYER M4 ;
      RECT 524.85 0.0 524.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[71]
  PIN QA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 52.19 0.0 52.33 0.39 ;
      LAYER M3 ;
      RECT 52.19 0.0 52.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[8]
  PIN DYA[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 525.62 0.0 525.76 0.39 ;
      LAYER M2 ;
      RECT 525.62 0.0 525.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[71]
  PIN DYA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 51.42 0.0 51.56 0.39 ;
      LAYER M1 ;
      RECT 51.42 0.0 51.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[8]
  PIN TDA[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 526.115 0.0 526.255 0.39 ;
      LAYER M4 ;
      RECT 526.115 0.0 526.255 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[71]
  PIN TDA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 50.925 0.0 51.065 0.39 ;
      LAYER M3 ;
      RECT 50.925 0.0 51.065 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[8]
  PIN TQA[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 526.4 0.0 526.54 0.39 ;
      LAYER M4 ;
      RECT 526.4 0.0 526.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[71]
  PIN TQA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 50.64 0.0 50.78 0.39 ;
      LAYER M3 ;
      RECT 50.64 0.0 50.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[8]
  PIN TQB[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 526.99 0.0 527.13 0.39 ;
      LAYER M4 ;
      RECT 526.99 0.0 527.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[72]
  PIN TQB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 50.05 0.0 50.19 0.39 ;
      LAYER M3 ;
      RECT 50.05 0.0 50.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[7]
  PIN TDB[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 527.24 0.0 527.38 0.39 ;
      LAYER M4 ;
      RECT 527.24 0.0 527.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[72]
  PIN TDB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 49.8 0.0 49.94 0.39 ;
      LAYER M3 ;
      RECT 49.8 0.0 49.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[7]
  PIN DYB[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 527.73 0.0 527.87 0.39 ;
      LAYER M2 ;
      RECT 527.73 0.0 527.87 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[72]
  PIN DYB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 49.31 0.0 49.45 0.39 ;
      LAYER M1 ;
      RECT 49.31 0.0 49.45 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[7]
  PIN QB[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 528.5 0.0 528.64 0.39 ;
      LAYER M4 ;
      RECT 528.5 0.0 528.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[72]
  PIN QB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 48.54 0.0 48.68 0.39 ;
      LAYER M3 ;
      RECT 48.54 0.0 48.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[7]
  PIN DB[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 529.49 0.0 529.63 0.39 ;
      LAYER M4 ;
      RECT 529.49 0.0 529.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[72]
  PIN DB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 47.55 0.0 47.69 0.39 ;
      LAYER M3 ;
      RECT 47.55 0.0 47.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[7]
  PIN DA[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 530.06 0.0 530.2 0.39 ;
      LAYER M4 ;
      RECT 530.06 0.0 530.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[72]
  PIN DA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 46.98 0.0 47.12 0.39 ;
      LAYER M3 ;
      RECT 46.98 0.0 47.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[7]
  PIN QA[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 531.05 0.0 531.19 0.39 ;
      LAYER M4 ;
      RECT 531.05 0.0 531.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[72]
  PIN QA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 45.99 0.0 46.13 0.39 ;
      LAYER M3 ;
      RECT 45.99 0.0 46.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[7]
  PIN DYA[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 531.82 0.0 531.96 0.39 ;
      LAYER M2 ;
      RECT 531.82 0.0 531.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[72]
  PIN DYA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 45.22 0.0 45.36 0.39 ;
      LAYER M1 ;
      RECT 45.22 0.0 45.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[7]
  PIN TDA[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 532.315 0.0 532.455 0.39 ;
      LAYER M4 ;
      RECT 532.315 0.0 532.455 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[72]
  PIN TDA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 44.725 0.0 44.865 0.39 ;
      LAYER M3 ;
      RECT 44.725 0.0 44.865 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[7]
  PIN TQA[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 532.6 0.0 532.74 0.39 ;
      LAYER M4 ;
      RECT 532.6 0.0 532.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[72]
  PIN TQA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 44.44 0.0 44.58 0.39 ;
      LAYER M3 ;
      RECT 44.44 0.0 44.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[7]
  PIN TQB[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 533.19 0.0 533.33 0.39 ;
      LAYER M4 ;
      RECT 533.19 0.0 533.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[73]
  PIN TQB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 43.85 0.0 43.99 0.39 ;
      LAYER M3 ;
      RECT 43.85 0.0 43.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[6]
  PIN TDB[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 533.44 0.0 533.58 0.39 ;
      LAYER M4 ;
      RECT 533.44 0.0 533.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[73]
  PIN TDB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 43.6 0.0 43.74 0.39 ;
      LAYER M3 ;
      RECT 43.6 0.0 43.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[6]
  PIN DYB[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 533.93 0.0 534.07 0.39 ;
      LAYER M2 ;
      RECT 533.93 0.0 534.07 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[73]
  PIN DYB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 43.11 0.0 43.25 0.39 ;
      LAYER M1 ;
      RECT 43.11 0.0 43.25 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[6]
  PIN QB[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 534.7 0.0 534.84 0.39 ;
      LAYER M4 ;
      RECT 534.7 0.0 534.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[73]
  PIN QB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 42.34 0.0 42.48 0.39 ;
      LAYER M3 ;
      RECT 42.34 0.0 42.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[6]
  PIN DB[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 535.69 0.0 535.83 0.39 ;
      LAYER M4 ;
      RECT 535.69 0.0 535.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[73]
  PIN DB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 41.35 0.0 41.49 0.39 ;
      LAYER M3 ;
      RECT 41.35 0.0 41.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[6]
  PIN DA[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 536.26 0.0 536.4 0.39 ;
      LAYER M4 ;
      RECT 536.26 0.0 536.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[73]
  PIN DA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 40.78 0.0 40.92 0.39 ;
      LAYER M3 ;
      RECT 40.78 0.0 40.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[6]
  PIN QA[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 537.25 0.0 537.39 0.39 ;
      LAYER M4 ;
      RECT 537.25 0.0 537.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[73]
  PIN QA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 39.79 0.0 39.93 0.39 ;
      LAYER M3 ;
      RECT 39.79 0.0 39.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[6]
  PIN DYA[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 538.02 0.0 538.16 0.39 ;
      LAYER M2 ;
      RECT 538.02 0.0 538.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[73]
  PIN DYA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 39.02 0.0 39.16 0.39 ;
      LAYER M1 ;
      RECT 39.02 0.0 39.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[6]
  PIN TDA[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 538.515 0.0 538.655 0.39 ;
      LAYER M4 ;
      RECT 538.515 0.0 538.655 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[73]
  PIN TDA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 38.525 0.0 38.665 0.39 ;
      LAYER M3 ;
      RECT 38.525 0.0 38.665 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[6]
  PIN TQA[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 538.8 0.0 538.94 0.39 ;
      LAYER M4 ;
      RECT 538.8 0.0 538.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[73]
  PIN TQA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 38.24 0.0 38.38 0.39 ;
      LAYER M3 ;
      RECT 38.24 0.0 38.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[6]
  PIN TQB[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 539.39 0.0 539.53 0.39 ;
      LAYER M4 ;
      RECT 539.39 0.0 539.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[74]
  PIN TQB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 37.65 0.0 37.79 0.39 ;
      LAYER M3 ;
      RECT 37.65 0.0 37.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[5]
  PIN TDB[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 539.64 0.0 539.78 0.39 ;
      LAYER M4 ;
      RECT 539.64 0.0 539.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[74]
  PIN TDB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 37.4 0.0 37.54 0.39 ;
      LAYER M3 ;
      RECT 37.4 0.0 37.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[5]
  PIN DYB[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 540.13 0.0 540.27 0.39 ;
      LAYER M2 ;
      RECT 540.13 0.0 540.27 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[74]
  PIN DYB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 36.91 0.0 37.05 0.39 ;
      LAYER M1 ;
      RECT 36.91 0.0 37.05 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[5]
  PIN QB[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 540.9 0.0 541.04 0.39 ;
      LAYER M4 ;
      RECT 540.9 0.0 541.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[74]
  PIN QB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 36.14 0.0 36.28 0.39 ;
      LAYER M3 ;
      RECT 36.14 0.0 36.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[5]
  PIN DB[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 541.89 0.0 542.03 0.39 ;
      LAYER M4 ;
      RECT 541.89 0.0 542.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[74]
  PIN DB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 35.15 0.0 35.29 0.39 ;
      LAYER M3 ;
      RECT 35.15 0.0 35.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[5]
  PIN DA[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 542.46 0.0 542.6 0.39 ;
      LAYER M4 ;
      RECT 542.46 0.0 542.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[74]
  PIN DA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 34.58 0.0 34.72 0.39 ;
      LAYER M3 ;
      RECT 34.58 0.0 34.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[5]
  PIN QA[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 543.45 0.0 543.59 0.39 ;
      LAYER M4 ;
      RECT 543.45 0.0 543.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[74]
  PIN QA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 33.59 0.0 33.73 0.39 ;
      LAYER M3 ;
      RECT 33.59 0.0 33.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[5]
  PIN DYA[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 544.22 0.0 544.36 0.39 ;
      LAYER M2 ;
      RECT 544.22 0.0 544.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[74]
  PIN DYA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 32.82 0.0 32.96 0.39 ;
      LAYER M1 ;
      RECT 32.82 0.0 32.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[5]
  PIN TDA[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 544.715 0.0 544.855 0.39 ;
      LAYER M4 ;
      RECT 544.715 0.0 544.855 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[74]
  PIN TDA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 32.325 0.0 32.465 0.39 ;
      LAYER M3 ;
      RECT 32.325 0.0 32.465 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[5]
  PIN TQA[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 545.0 0.0 545.14 0.39 ;
      LAYER M4 ;
      RECT 545.0 0.0 545.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[74]
  PIN TQA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 32.04 0.0 32.18 0.39 ;
      LAYER M3 ;
      RECT 32.04 0.0 32.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[5]
  PIN TQB[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 545.59 0.0 545.73 0.39 ;
      LAYER M4 ;
      RECT 545.59 0.0 545.73 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[75]
  PIN TQB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 31.45 0.0 31.59 0.39 ;
      LAYER M3 ;
      RECT 31.45 0.0 31.59 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[4]
  PIN TDB[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 545.84 0.0 545.98 0.39 ;
      LAYER M4 ;
      RECT 545.84 0.0 545.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[75]
  PIN TDB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 31.2 0.0 31.34 0.39 ;
      LAYER M3 ;
      RECT 31.2 0.0 31.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[4]
  PIN DYB[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 546.33 0.0 546.47 0.39 ;
      LAYER M2 ;
      RECT 546.33 0.0 546.47 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[75]
  PIN DYB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 30.71 0.0 30.85 0.39 ;
      LAYER M1 ;
      RECT 30.71 0.0 30.85 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[4]
  PIN QB[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 547.1 0.0 547.24 0.39 ;
      LAYER M4 ;
      RECT 547.1 0.0 547.24 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[75]
  PIN QB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 29.94 0.0 30.08 0.39 ;
      LAYER M3 ;
      RECT 29.94 0.0 30.08 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[4]
  PIN DB[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 548.09 0.0 548.23 0.39 ;
      LAYER M4 ;
      RECT 548.09 0.0 548.23 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[75]
  PIN DB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 28.95 0.0 29.09 0.39 ;
      LAYER M3 ;
      RECT 28.95 0.0 29.09 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[4]
  PIN DA[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 548.66 0.0 548.8 0.39 ;
      LAYER M4 ;
      RECT 548.66 0.0 548.8 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[75]
  PIN DA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 28.38 0.0 28.52 0.39 ;
      LAYER M3 ;
      RECT 28.38 0.0 28.52 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[4]
  PIN QA[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 549.65 0.0 549.79 0.39 ;
      LAYER M4 ;
      RECT 549.65 0.0 549.79 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[75]
  PIN QA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 27.39 0.0 27.53 0.39 ;
      LAYER M3 ;
      RECT 27.39 0.0 27.53 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[4]
  PIN DYA[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 550.42 0.0 550.56 0.39 ;
      LAYER M2 ;
      RECT 550.42 0.0 550.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[75]
  PIN DYA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 26.62 0.0 26.76 0.39 ;
      LAYER M1 ;
      RECT 26.62 0.0 26.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[4]
  PIN TDA[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 550.915 0.0 551.055 0.39 ;
      LAYER M4 ;
      RECT 550.915 0.0 551.055 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[75]
  PIN TDA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 26.125 0.0 26.265 0.39 ;
      LAYER M3 ;
      RECT 26.125 0.0 26.265 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[4]
  PIN TQA[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 551.2 0.0 551.34 0.39 ;
      LAYER M4 ;
      RECT 551.2 0.0 551.34 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[75]
  PIN TQA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 25.84 0.0 25.98 0.39 ;
      LAYER M3 ;
      RECT 25.84 0.0 25.98 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[4]
  PIN TQB[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 551.79 0.0 551.93 0.39 ;
      LAYER M4 ;
      RECT 551.79 0.0 551.93 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[76]
  PIN TQB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 25.25 0.0 25.39 0.39 ;
      LAYER M3 ;
      RECT 25.25 0.0 25.39 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[3]
  PIN TDB[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 552.04 0.0 552.18 0.39 ;
      LAYER M4 ;
      RECT 552.04 0.0 552.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[76]
  PIN TDB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 25.0 0.0 25.14 0.39 ;
      LAYER M3 ;
      RECT 25.0 0.0 25.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[3]
  PIN DYB[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 552.53 0.0 552.67 0.39 ;
      LAYER M2 ;
      RECT 552.53 0.0 552.67 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[76]
  PIN DYB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 24.51 0.0 24.65 0.39 ;
      LAYER M1 ;
      RECT 24.51 0.0 24.65 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[3]
  PIN QB[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 553.3 0.0 553.44 0.39 ;
      LAYER M4 ;
      RECT 553.3 0.0 553.44 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[76]
  PIN QB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 23.74 0.0 23.88 0.39 ;
      LAYER M3 ;
      RECT 23.74 0.0 23.88 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[3]
  PIN DB[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 554.29 0.0 554.43 0.39 ;
      LAYER M4 ;
      RECT 554.29 0.0 554.43 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[76]
  PIN DB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 22.75 0.0 22.89 0.39 ;
      LAYER M3 ;
      RECT 22.75 0.0 22.89 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[3]
  PIN DA[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 554.86 0.0 555.0 0.39 ;
      LAYER M4 ;
      RECT 554.86 0.0 555.0 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[76]
  PIN DA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 22.18 0.0 22.32 0.39 ;
      LAYER M3 ;
      RECT 22.18 0.0 22.32 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[3]
  PIN QA[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 555.85 0.0 555.99 0.39 ;
      LAYER M4 ;
      RECT 555.85 0.0 555.99 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[76]
  PIN QA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 21.19 0.0 21.33 0.39 ;
      LAYER M3 ;
      RECT 21.19 0.0 21.33 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[3]
  PIN DYA[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 556.62 0.0 556.76 0.39 ;
      LAYER M2 ;
      RECT 556.62 0.0 556.76 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[76]
  PIN DYA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 20.42 0.0 20.56 0.39 ;
      LAYER M1 ;
      RECT 20.42 0.0 20.56 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[3]
  PIN TDA[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 557.115 0.0 557.255 0.39 ;
      LAYER M4 ;
      RECT 557.115 0.0 557.255 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[76]
  PIN TDA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 19.925 0.0 20.065 0.39 ;
      LAYER M3 ;
      RECT 19.925 0.0 20.065 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[3]
  PIN TQA[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 557.4 0.0 557.54 0.39 ;
      LAYER M4 ;
      RECT 557.4 0.0 557.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[76]
  PIN TQA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 19.64 0.0 19.78 0.39 ;
      LAYER M3 ;
      RECT 19.64 0.0 19.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[3]
  PIN TQB[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 557.99 0.0 558.13 0.39 ;
      LAYER M4 ;
      RECT 557.99 0.0 558.13 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[77]
  PIN TQB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 19.05 0.0 19.19 0.39 ;
      LAYER M3 ;
      RECT 19.05 0.0 19.19 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[2]
  PIN TDB[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 558.24 0.0 558.38 0.39 ;
      LAYER M4 ;
      RECT 558.24 0.0 558.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[77]
  PIN TDB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 18.8 0.0 18.94 0.39 ;
      LAYER M3 ;
      RECT 18.8 0.0 18.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[2]
  PIN DYB[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 558.73 0.0 558.87 0.39 ;
      LAYER M2 ;
      RECT 558.73 0.0 558.87 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[77]
  PIN DYB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 18.31 0.0 18.45 0.39 ;
      LAYER M1 ;
      RECT 18.31 0.0 18.45 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[2]
  PIN QB[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 559.5 0.0 559.64 0.39 ;
      LAYER M4 ;
      RECT 559.5 0.0 559.64 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[77]
  PIN QB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 17.54 0.0 17.68 0.39 ;
      LAYER M3 ;
      RECT 17.54 0.0 17.68 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[2]
  PIN DB[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 560.49 0.0 560.63 0.39 ;
      LAYER M4 ;
      RECT 560.49 0.0 560.63 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[77]
  PIN DB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 16.55 0.0 16.69 0.39 ;
      LAYER M3 ;
      RECT 16.55 0.0 16.69 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[2]
  PIN DA[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 561.06 0.0 561.2 0.39 ;
      LAYER M4 ;
      RECT 561.06 0.0 561.2 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[77]
  PIN DA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 15.98 0.0 16.12 0.39 ;
      LAYER M3 ;
      RECT 15.98 0.0 16.12 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[2]
  PIN QA[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 562.05 0.0 562.19 0.39 ;
      LAYER M4 ;
      RECT 562.05 0.0 562.19 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[77]
  PIN QA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 14.99 0.0 15.13 0.39 ;
      LAYER M3 ;
      RECT 14.99 0.0 15.13 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[2]
  PIN DYA[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 562.82 0.0 562.96 0.39 ;
      LAYER M2 ;
      RECT 562.82 0.0 562.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[77]
  PIN DYA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 14.22 0.0 14.36 0.39 ;
      LAYER M1 ;
      RECT 14.22 0.0 14.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[2]
  PIN TDA[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 563.315 0.0 563.455 0.39 ;
      LAYER M4 ;
      RECT 563.315 0.0 563.455 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[77]
  PIN TDA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 13.725 0.0 13.865 0.39 ;
      LAYER M3 ;
      RECT 13.725 0.0 13.865 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[2]
  PIN TQA[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 563.6 0.0 563.74 0.39 ;
      LAYER M4 ;
      RECT 563.6 0.0 563.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[77]
  PIN TQA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 13.44 0.0 13.58 0.39 ;
      LAYER M3 ;
      RECT 13.44 0.0 13.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[2]
  PIN TQB[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 564.19 0.0 564.33 0.39 ;
      LAYER M4 ;
      RECT 564.19 0.0 564.33 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[78]
  PIN TQB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 12.85 0.0 12.99 0.39 ;
      LAYER M3 ;
      RECT 12.85 0.0 12.99 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[1]
  PIN TDB[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 564.44 0.0 564.58 0.39 ;
      LAYER M4 ;
      RECT 564.44 0.0 564.58 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[78]
  PIN TDB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 12.6 0.0 12.74 0.39 ;
      LAYER M3 ;
      RECT 12.6 0.0 12.74 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[1]
  PIN DYB[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 564.93 0.0 565.07 0.39 ;
      LAYER M2 ;
      RECT 564.93 0.0 565.07 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[78]
  PIN DYB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 12.11 0.0 12.25 0.39 ;
      LAYER M1 ;
      RECT 12.11 0.0 12.25 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[1]
  PIN QB[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 565.7 0.0 565.84 0.39 ;
      LAYER M4 ;
      RECT 565.7 0.0 565.84 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[78]
  PIN QB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.34 0.0 11.48 0.39 ;
      LAYER M3 ;
      RECT 11.34 0.0 11.48 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[1]
  PIN DB[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 566.69 0.0 566.83 0.39 ;
      LAYER M4 ;
      RECT 566.69 0.0 566.83 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[78]
  PIN DB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.35 0.0 10.49 0.39 ;
      LAYER M3 ;
      RECT 10.35 0.0 10.49 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[1]
  PIN DA[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 567.26 0.0 567.4 0.39 ;
      LAYER M4 ;
      RECT 567.26 0.0 567.4 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[78]
  PIN DA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 9.78 0.0 9.92 0.39 ;
      LAYER M3 ;
      RECT 9.78 0.0 9.92 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[1]
  PIN QA[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 568.25 0.0 568.39 0.39 ;
      LAYER M4 ;
      RECT 568.25 0.0 568.39 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[78]
  PIN QA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 8.79 0.0 8.93 0.39 ;
      LAYER M3 ;
      RECT 8.79 0.0 8.93 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[1]
  PIN DYA[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 569.02 0.0 569.16 0.39 ;
      LAYER M2 ;
      RECT 569.02 0.0 569.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[78]
  PIN DYA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 8.02 0.0 8.16 0.39 ;
      LAYER M1 ;
      RECT 8.02 0.0 8.16 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[1]
  PIN TDA[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 569.515 0.0 569.655 0.39 ;
      LAYER M4 ;
      RECT 569.515 0.0 569.655 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[78]
  PIN TDA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 7.525 0.0 7.665 0.39 ;
      LAYER M3 ;
      RECT 7.525 0.0 7.665 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[1]
  PIN TQA[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 569.8 0.0 569.94 0.39 ;
      LAYER M4 ;
      RECT 569.8 0.0 569.94 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[78]
  PIN TQA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 7.24 0.0 7.38 0.39 ;
      LAYER M3 ;
      RECT 7.24 0.0 7.38 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[1]
  PIN TQB[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 570.39 0.0 570.53 0.39 ;
      LAYER M4 ;
      RECT 570.39 0.0 570.53 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[79]
  PIN TQB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 6.65 0.0 6.79 0.39 ;
      LAYER M3 ;
      RECT 6.65 0.0 6.79 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQB[0]
  PIN TDB[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 570.64 0.0 570.78 0.39 ;
      LAYER M4 ;
      RECT 570.64 0.0 570.78 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[79]
  PIN TDB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 6.4 0.0 6.54 0.39 ;
      LAYER M3 ;
      RECT 6.4 0.0 6.54 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDB[0]
  PIN DYB[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 571.13 0.0 571.27 0.39 ;
      LAYER M2 ;
      RECT 571.13 0.0 571.27 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[79]
  PIN DYB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 5.91 0.0 6.05 0.39 ;
      LAYER M1 ;
      RECT 5.91 0.0 6.05 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYB[0]
  PIN QB[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 571.9 0.0 572.04 0.39 ;
      LAYER M4 ;
      RECT 571.9 0.0 572.04 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[79]
  PIN QB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 5.14 0.0 5.28 0.39 ;
      LAYER M3 ;
      RECT 5.14 0.0 5.28 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QB[0]
  PIN DB[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 572.89 0.0 573.03 0.39 ;
      LAYER M4 ;
      RECT 572.89 0.0 573.03 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[79]
  PIN DB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 4.15 0.0 4.29 0.39 ;
      LAYER M3 ;
      RECT 4.15 0.0 4.29 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DB[0]
  PIN DA[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 573.46 0.0 573.6 0.39 ;
      LAYER M4 ;
      RECT 573.46 0.0 573.6 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[79]
  PIN DA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 3.58 0.0 3.72 0.39 ;
      LAYER M3 ;
      RECT 3.58 0.0 3.72 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END DA[0]
  PIN QA[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 574.45 0.0 574.59 0.39 ;
      LAYER M4 ;
      RECT 574.45 0.0 574.59 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[79]
  PIN QA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 2.59 0.0 2.73 0.39 ;
      LAYER M3 ;
      RECT 2.59 0.0 2.73 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END QA[0]
  PIN DYA[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 575.22 0.0 575.36 0.39 ;
      LAYER M2 ;
      RECT 575.22 0.0 575.36 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[79]
  PIN DYA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 1.82 0.0 1.96 0.39 ;
      LAYER M1 ;
      RECT 1.82 0.0 1.96 0.39 ;
      END
    ANTENNADIFFAREA 0.06 ;
    END DYA[0]
  PIN TDA[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 575.715 0.0 575.855 0.39 ;
      LAYER M4 ;
      RECT 575.715 0.0 575.855 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[79]
  PIN TDA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 1.325 0.0 1.465 0.39 ;
      LAYER M3 ;
      RECT 1.325 0.0 1.465 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TDA[0]
  PIN TQA[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 576.0 0.0 576.14 0.39 ;
      LAYER M4 ;
      RECT 576.0 0.0 576.14 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[79]
  PIN TQA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 1.04 0.0 1.18 0.39 ;
      LAYER M3 ;
      RECT 1.04 0.0 1.18 0.39 ;
      END
    ANTENNAGATEAREA 0.009 ;
    ANTENNADIFFAREA 0.06 ;
    END TQA[0]
  PIN VDDCE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 3.83 0.0 4.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.03 0.0 10.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 16.23 0.0 16.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 22.43 0.0 22.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.63 0.0 28.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 34.83 0.0 35.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 41.03 0.0 41.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.23 0.0 47.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 53.43 0.0 53.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 59.63 0.0 59.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 65.83 0.0 66.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.03 0.0 72.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.23 0.0 78.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.43 0.0 84.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.63 0.0 90.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 96.83 0.0 97.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.03 0.0 103.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 109.23 0.0 109.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 115.43 0.0 115.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 121.63 0.0 121.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 126.065 0.0 126.275 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 129.4 0.0 129.61 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 134.045 0.0 134.255 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 137.505 0.0 137.715 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 140.795 0.0 141.005 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.875 0.0 148.085 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 151.165 0.0 151.375 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 154.625 0.0 154.835 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 159.27 0.0 159.48 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 162.605 0.0 162.815 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 167.04 0.0 167.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 173.24 0.0 173.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 179.44 0.0 179.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 185.64 0.0 185.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 191.84 0.0 192.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 198.04 0.0 198.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 204.24 0.0 204.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 210.44 0.0 210.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 216.64 0.0 216.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 222.84 0.0 223.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.04 0.0 229.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.24 0.0 235.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 241.44 0.0 241.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 247.64 0.0 247.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 253.84 0.0 254.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 260.04 0.0 260.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 266.24 0.0 266.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 272.44 0.0 272.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 278.64 0.0 278.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 284.84 0.0 285.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 292.13 0.0 292.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 298.33 0.0 298.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 304.53 0.0 304.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 310.73 0.0 310.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 316.93 0.0 317.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 323.13 0.0 323.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 329.33 0.0 329.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 335.53 0.0 335.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 341.73 0.0 341.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 347.93 0.0 348.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 354.13 0.0 354.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 360.33 0.0 360.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 366.53 0.0 366.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 372.73 0.0 372.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 378.93 0.0 379.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 385.13 0.0 385.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 391.33 0.0 391.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 397.53 0.0 397.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 403.73 0.0 403.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 409.93 0.0 410.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 414.365 0.0 414.575 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 417.7 0.0 417.91 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 422.345 0.0 422.555 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 425.805 0.0 426.015 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 429.095 0.0 429.305 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 436.175 0.0 436.385 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 439.465 0.0 439.675 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 442.925 0.0 443.135 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 447.57 0.0 447.78 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 450.905 0.0 451.115 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 455.34 0.0 455.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 461.54 0.0 461.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 467.74 0.0 467.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 473.94 0.0 474.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 480.14 0.0 480.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 486.34 0.0 486.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 492.54 0.0 492.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 498.74 0.0 498.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 504.94 0.0 505.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 511.14 0.0 511.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 517.34 0.0 517.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 523.54 0.0 523.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 529.74 0.0 529.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 535.94 0.0 536.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 542.14 0.0 542.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 548.34 0.0 548.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 554.54 0.0 554.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 560.74 0.0 560.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 566.94 0.0 567.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 573.14 0.0 573.35 270.08 ;
      END
    END VDDCE
  PIN VDDPE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.38 0.0 0.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 1.57 0.0 1.78 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 6.09 0.0 6.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.77 0.0 7.98 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.29 0.0 12.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 13.97 0.0 14.18 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 18.49 0.0 18.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.17 0.0 20.38 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 24.69 0.0 24.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 26.37 0.0 26.58 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.89 0.0 31.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.57 0.0 32.78 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.09 0.0 37.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.77 0.0 38.98 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 43.29 0.0 43.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.97 0.0 45.18 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 49.49 0.0 49.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.17 0.0 51.38 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.69 0.0 55.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 57.37 0.0 57.58 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.89 0.0 62.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 63.57 0.0 63.78 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.09 0.0 68.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 69.77 0.0 69.98 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.29 0.0 74.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.97 0.0 76.18 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 80.49 0.0 80.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.17 0.0 82.38 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 86.69 0.0 86.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.37 0.0 88.58 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.89 0.0 93.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.57 0.0 94.78 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 99.09 0.0 99.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.77 0.0 100.98 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 105.29 0.0 105.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 106.97 0.0 107.18 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 111.49 0.0 111.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 113.17 0.0 113.38 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 117.69 0.0 117.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 119.37 0.0 119.58 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.89 0.0 124.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.335 0.0 128.545 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 132.06 0.0 132.27 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 136.17 0.0 136.66 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 139.415 0.0 139.625 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 141.705 0.0 141.915 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 146.965 0.0 147.175 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 149.255 0.0 149.465 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 152.5 0.0 152.71 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.61 0.0 156.82 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 160.335 0.0 160.545 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 164.78 0.0 164.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 169.3 0.0 169.51 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 170.98 0.0 171.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 175.5 0.0 175.71 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.18 0.0 177.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 181.7 0.0 181.91 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 183.38 0.0 183.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.9 0.0 188.11 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 189.58 0.0 189.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 194.1 0.0 194.31 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 195.78 0.0 195.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 200.3 0.0 200.51 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 201.98 0.0 202.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 206.5 0.0 206.71 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 208.18 0.0 208.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 212.7 0.0 212.91 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 214.38 0.0 214.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 218.9 0.0 219.11 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 220.58 0.0 220.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.1 0.0 225.31 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 226.78 0.0 226.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 231.3 0.0 231.51 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.98 0.0 233.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 237.5 0.0 237.71 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.18 0.0 239.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 243.7 0.0 243.91 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 245.38 0.0 245.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.9 0.0 250.11 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 251.58 0.0 251.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 256.1 0.0 256.31 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 257.78 0.0 257.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.3 0.0 262.51 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 263.98 0.0 264.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 268.5 0.0 268.71 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 270.18 0.0 270.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 274.7 0.0 274.91 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 276.38 0.0 276.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 280.9 0.0 281.11 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 282.58 0.0 282.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 287.1 0.0 287.31 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 289.87 0.0 290.08 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 294.39 0.0 294.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 296.07 0.0 296.28 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 300.59 0.0 300.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 302.27 0.0 302.48 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 306.79 0.0 307.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 308.47 0.0 308.68 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 312.99 0.0 313.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 314.67 0.0 314.88 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 319.19 0.0 319.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 320.87 0.0 321.08 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 325.39 0.0 325.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 327.07 0.0 327.28 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 331.59 0.0 331.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 333.27 0.0 333.48 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 337.79 0.0 338.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 339.47 0.0 339.68 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 343.99 0.0 344.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 345.67 0.0 345.88 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 350.19 0.0 350.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 351.87 0.0 352.08 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 356.39 0.0 356.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 358.07 0.0 358.28 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 362.59 0.0 362.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 364.27 0.0 364.48 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 368.79 0.0 369.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 370.47 0.0 370.68 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 374.99 0.0 375.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 376.67 0.0 376.88 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 381.19 0.0 381.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 382.87 0.0 383.08 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 387.39 0.0 387.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 389.07 0.0 389.28 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 393.59 0.0 393.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 395.27 0.0 395.48 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 399.79 0.0 400.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 401.47 0.0 401.68 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 405.99 0.0 406.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 407.67 0.0 407.88 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 412.19 0.0 412.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 416.635 0.0 416.845 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 420.36 0.0 420.57 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 424.47 0.0 424.68 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 427.715 0.0 427.925 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 430.005 0.0 430.215 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 435.265 0.0 435.475 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 437.555 0.0 437.765 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 440.52 0.0 441.01 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 444.91 0.0 445.12 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 448.635 0.0 448.845 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 453.08 0.0 453.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 457.6 0.0 457.81 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 459.28 0.0 459.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 463.8 0.0 464.01 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 465.48 0.0 465.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 470.0 0.0 470.21 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 471.68 0.0 471.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 476.2 0.0 476.41 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 477.88 0.0 478.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 482.4 0.0 482.61 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 484.08 0.0 484.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 488.6 0.0 488.81 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 490.28 0.0 490.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 494.8 0.0 495.01 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 496.48 0.0 496.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 501.0 0.0 501.21 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 502.68 0.0 502.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 507.2 0.0 507.41 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 508.88 0.0 509.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 513.4 0.0 513.61 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 515.08 0.0 515.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 519.6 0.0 519.81 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 521.28 0.0 521.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 525.8 0.0 526.01 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 527.48 0.0 527.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 532.0 0.0 532.21 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 533.68 0.0 533.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 538.2 0.0 538.41 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 539.88 0.0 540.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 544.4 0.0 544.61 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 546.08 0.0 546.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 550.6 0.0 550.81 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 552.28 0.0 552.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 556.8 0.0 557.01 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 558.48 0.0 558.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 563.0 0.0 563.21 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 564.68 0.0 564.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 569.2 0.0 569.41 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 570.88 0.0 571.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 575.4 0.0 575.61 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 576.59 0.0 576.8 270.08 ;
      END
    END VDDPE
  PIN VSSE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.73 0.0 0.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 2.28 0.0 2.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 5.38 0.0 5.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 6.93 0.0 7.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 8.48 0.0 8.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 11.58 0.0 11.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 13.13 0.0 13.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 14.68 0.0 14.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.78 0.0 17.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.33 0.0 19.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.88 0.0 21.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 23.98 0.0 24.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.53 0.0 25.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.08 0.0 27.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.18 0.0 30.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 31.73 0.0 31.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 33.28 0.0 33.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 36.38 0.0 36.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.93 0.0 38.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 39.48 0.0 39.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.58 0.0 42.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.13 0.0 44.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.68 0.0 45.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.78 0.0 48.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.33 0.0 50.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.88 0.0 52.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 54.98 0.0 55.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 56.53 0.0 56.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.08 0.0 58.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.18 0.0 61.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 62.73 0.0 62.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.28 0.0 64.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.38 0.0 67.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.93 0.0 69.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.48 0.0 70.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 73.58 0.0 73.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.13 0.0 75.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 76.68 0.0 76.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 79.78 0.0 79.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.33 0.0 81.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.88 0.0 83.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 85.98 0.0 86.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.53 0.0 87.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 89.08 0.0 89.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.18 0.0 92.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 93.73 0.0 93.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 95.28 0.0 95.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.38 0.0 98.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 99.93 0.0 100.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 101.48 0.0 101.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 104.58 0.0 104.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 106.13 0.0 106.34 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 107.68 0.0 107.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 110.78 0.0 110.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 112.33 0.0 112.54 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 113.88 0.0 114.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 116.98 0.0 117.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.53 0.0 118.74 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.08 0.0 120.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.18 0.0 123.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 124.73 0.0 124.94 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 126.455 0.0 126.665 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 132.38 0.0 132.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 134.365 0.0 134.575 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 137.825 0.0 138.035 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 138.525 0.0 138.735 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 140.475 0.0 140.685 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.74 0.0 143.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.93 0.0 145.14 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 148.195 0.0 148.405 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 150.145 0.0 150.355 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 150.845 0.0 151.055 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 154.305 0.0 154.515 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.29 0.0 156.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 162.215 0.0 162.425 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 163.94 0.0 164.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 165.49 0.0 165.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 168.59 0.0 168.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 170.14 0.0 170.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 171.69 0.0 171.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 174.79 0.0 175.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 176.34 0.0 176.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.89 0.0 178.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 180.99 0.0 181.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 182.54 0.0 182.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 184.09 0.0 184.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.19 0.0 187.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 188.74 0.0 188.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.29 0.0 190.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 193.39 0.0 193.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 194.94 0.0 195.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.49 0.0 196.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.59 0.0 199.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 201.14 0.0 201.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 202.69 0.0 202.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 205.79 0.0 206.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.34 0.0 207.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 208.89 0.0 209.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 211.99 0.0 212.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.54 0.0 213.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.09 0.0 215.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 218.19 0.0 218.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 219.74 0.0 219.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 221.29 0.0 221.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 224.39 0.0 224.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.94 0.0 226.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 227.49 0.0 227.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 230.59 0.0 230.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.14 0.0 232.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 233.69 0.0 233.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 236.79 0.0 237.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 238.34 0.0 238.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.89 0.0 240.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.99 0.0 243.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 244.54 0.0 244.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 246.09 0.0 246.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.19 0.0 249.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 250.74 0.0 250.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.29 0.0 252.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 255.39 0.0 255.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 256.94 0.0 257.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 258.49 0.0 258.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 261.59 0.0 261.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 263.14 0.0 263.35 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 264.69 0.0 264.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 267.79 0.0 268.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 269.34 0.0 269.55 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 270.89 0.0 271.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 273.99 0.0 274.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 275.54 0.0 275.75 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 277.09 0.0 277.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 280.19 0.0 280.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 281.74 0.0 281.95 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 283.29 0.0 283.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 286.39 0.0 286.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 287.94 0.0 288.15 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 289.03 0.0 289.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 290.58 0.0 290.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 293.68 0.0 293.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 295.23 0.0 295.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 296.78 0.0 296.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 299.88 0.0 300.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 301.43 0.0 301.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 302.98 0.0 303.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 306.08 0.0 306.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 307.63 0.0 307.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 309.18 0.0 309.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 312.28 0.0 312.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 313.83 0.0 314.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 315.38 0.0 315.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 318.48 0.0 318.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 320.03 0.0 320.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 321.58 0.0 321.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 324.68 0.0 324.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 326.23 0.0 326.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 327.78 0.0 327.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 330.88 0.0 331.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 332.43 0.0 332.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 333.98 0.0 334.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 337.08 0.0 337.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 338.63 0.0 338.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 340.18 0.0 340.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 343.28 0.0 343.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 344.83 0.0 345.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 346.38 0.0 346.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 349.48 0.0 349.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 351.03 0.0 351.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 352.58 0.0 352.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 355.68 0.0 355.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 357.23 0.0 357.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 358.78 0.0 358.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 361.88 0.0 362.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 363.43 0.0 363.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 364.98 0.0 365.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 368.08 0.0 368.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 369.63 0.0 369.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 371.18 0.0 371.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 374.28 0.0 374.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 375.83 0.0 376.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 377.38 0.0 377.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 380.48 0.0 380.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 382.03 0.0 382.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 383.58 0.0 383.79 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 386.68 0.0 386.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 388.23 0.0 388.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 389.78 0.0 389.99 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 392.88 0.0 393.09 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 394.43 0.0 394.64 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 395.98 0.0 396.19 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 399.08 0.0 399.29 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 400.63 0.0 400.84 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 402.18 0.0 402.39 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 405.28 0.0 405.49 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 406.83 0.0 407.04 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 408.38 0.0 408.59 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 411.48 0.0 411.69 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 413.03 0.0 413.24 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 414.755 0.0 414.965 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 420.68 0.0 420.89 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 422.665 0.0 422.875 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 426.125 0.0 426.335 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 426.825 0.0 427.035 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 428.775 0.0 428.985 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 432.04 0.0 432.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 433.23 0.0 433.44 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 436.495 0.0 436.705 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 438.445 0.0 438.655 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 439.145 0.0 439.355 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 442.605 0.0 442.815 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 444.59 0.0 444.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 450.515 0.0 450.725 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 452.24 0.0 452.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 453.79 0.0 454.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 456.89 0.0 457.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 458.44 0.0 458.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 459.99 0.0 460.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 463.09 0.0 463.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 464.64 0.0 464.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 466.19 0.0 466.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 469.29 0.0 469.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 470.84 0.0 471.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 472.39 0.0 472.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 475.49 0.0 475.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 477.04 0.0 477.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 478.59 0.0 478.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 481.69 0.0 481.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 483.24 0.0 483.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 484.79 0.0 485.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 487.89 0.0 488.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 489.44 0.0 489.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 490.99 0.0 491.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 494.09 0.0 494.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 495.64 0.0 495.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 497.19 0.0 497.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 500.29 0.0 500.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 501.84 0.0 502.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 503.39 0.0 503.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 506.49 0.0 506.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 508.04 0.0 508.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 509.59 0.0 509.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 512.69 0.0 512.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 514.24 0.0 514.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 515.79 0.0 516.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 518.89 0.0 519.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 520.44 0.0 520.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 521.99 0.0 522.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 525.09 0.0 525.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 526.64 0.0 526.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 528.19 0.0 528.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 531.29 0.0 531.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 532.84 0.0 533.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 534.39 0.0 534.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 537.49 0.0 537.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 539.04 0.0 539.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 540.59 0.0 540.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 543.69 0.0 543.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 545.24 0.0 545.45 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 546.79 0.0 547.0 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 549.89 0.0 550.1 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 551.44 0.0 551.65 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 552.99 0.0 553.2 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 556.09 0.0 556.3 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 557.64 0.0 557.85 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 559.19 0.0 559.4 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 562.29 0.0 562.5 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 563.84 0.0 564.05 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 565.39 0.0 565.6 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 568.49 0.0 568.7 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 570.04 0.0 570.25 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 571.59 0.0 571.8 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 574.69 0.0 574.9 270.08 ;
      END
    PORT
      LAYER M4 ;
      RECT 576.24 0.0 576.45 270.08 ;
      END
    END VSSE
  OBS
    #otc obstructions
    LAYER M1 DESIGNRULEWIDTH 0.07 ;
    RECT 575.43 0.0 577.18 0.46 ;
    RECT 571.34 0.0 575.15 0.46 ;
    RECT 569.23 0.0 571.06 0.46 ;
    RECT 565.14 0.0 568.95 0.46 ;
    RECT 563.03 0.0 564.86 0.46 ;
    RECT 558.94 0.0 562.75 0.46 ;
    RECT 556.83 0.0 558.66 0.46 ;
    RECT 552.74 0.0 556.55 0.46 ;
    RECT 550.63 0.0 552.46 0.46 ;
    RECT 546.54 0.0 550.35 0.46 ;
    RECT 544.43 0.0 546.26 0.46 ;
    RECT 540.34 0.0 544.15 0.46 ;
    RECT 538.23 0.0 540.06 0.46 ;
    RECT 534.14 0.0 537.95 0.46 ;
    RECT 532.03 0.0 533.86 0.46 ;
    RECT 527.94 0.0 531.75 0.46 ;
    RECT 525.83 0.0 527.66 0.46 ;
    RECT 521.74 0.0 525.55 0.46 ;
    RECT 519.63 0.0 521.46 0.46 ;
    RECT 515.54 0.0 519.35 0.46 ;
    RECT 513.43 0.0 515.26 0.46 ;
    RECT 509.34 0.0 513.15 0.46 ;
    RECT 507.23 0.0 509.06 0.46 ;
    RECT 503.14 0.0 506.95 0.46 ;
    RECT 501.03 0.0 502.86 0.46 ;
    RECT 496.94 0.0 500.75 0.46 ;
    RECT 494.83 0.0 496.66 0.46 ;
    RECT 490.74 0.0 494.55 0.46 ;
    RECT 488.63 0.0 490.46 0.46 ;
    RECT 484.54 0.0 488.35 0.46 ;
    RECT 482.43 0.0 484.26 0.46 ;
    RECT 478.34 0.0 482.15 0.46 ;
    RECT 476.23 0.0 478.06 0.46 ;
    RECT 472.14 0.0 475.95 0.46 ;
    RECT 470.03 0.0 471.86 0.46 ;
    RECT 465.94 0.0 469.75 0.46 ;
    RECT 463.83 0.0 465.66 0.46 ;
    RECT 459.74 0.0 463.55 0.46 ;
    RECT 457.63 0.0 459.46 0.46 ;
    RECT 453.54 0.0 457.35 0.46 ;
    RECT 412.22 0.0 453.26 0.46 ;
    RECT 408.13 0.0 411.94 0.46 ;
    RECT 406.02 0.0 407.85 0.46 ;
    RECT 401.93 0.0 405.74 0.46 ;
    RECT 400.63 0.0 401.65 0.46 ;
    RECT 400.085 0.0 400.35 0.46 ;
    RECT 397.65 0.0 399.52 0.46 ;
    RECT 396.72 0.0 397.37 0.46 ;
    RECT 395.75 0.0 396.17 0.46 ;
    RECT 394.885 0.0 395.17 0.46 ;
    RECT 393.865 0.0 394.265 0.46 ;
    RECT 392.96 0.0 393.32 0.46 ;
    RECT 391.325 0.0 392.68 0.46 ;
    RECT 390.47 0.0 391.045 0.46 ;
    RECT 389.55 0.0 390.19 0.46 ;
    RECT 387.4 0.0 389.27 0.46 ;
    RECT 385.61 0.0 387.12 0.46 ;
    RECT 383.35 0.0 385.33 0.46 ;
    RECT 382.53 0.0 383.07 0.46 ;
    RECT 381.475 0.0 382.25 0.46 ;
    RECT 380.66 0.0 380.92 0.46 ;
    RECT 378.92 0.0 380.38 0.46 ;
    RECT 377.99 0.0 378.64 0.46 ;
    RECT 377.15 0.0 377.71 0.46 ;
    RECT 376.305 0.0 376.87 0.46 ;
    RECT 375.0 0.0 375.505 0.46 ;
    RECT 374.19 0.0 374.72 0.46 ;
    RECT 370.95 0.0 373.91 0.46 ;
    RECT 368.8 0.0 370.385 0.46 ;
    RECT 364.75 0.0 368.52 0.46 ;
    RECT 362.6 0.0 364.47 0.46 ;
    RECT 361.74 0.0 362.32 0.46 ;
    RECT 359.22 0.0 361.46 0.46 ;
    RECT 358.55 0.0 358.94 0.46 ;
    RECT 357.34 0.0 358.27 0.46 ;
    RECT 356.725 0.0 357.06 0.46 ;
    RECT 355.795 0.0 356.12 0.46 ;
    RECT 354.53 0.0 355.515 0.46 ;
    RECT 352.35 0.0 354.25 0.46 ;
    RECT 351.555 0.0 352.07 0.46 ;
    RECT 350.2 0.0 351.275 0.46 ;
    RECT 346.15 0.0 349.92 0.46 ;
    RECT 344.0 0.0 345.87 0.46 ;
    RECT 341.79 0.0 343.72 0.46 ;
    RECT 339.95 0.0 341.51 0.46 ;
    RECT 338.955 0.0 339.67 0.46 ;
    RECT 338.065 0.0 338.675 0.46 ;
    RECT 336.835 0.0 337.52 0.46 ;
    RECT 334.655 0.0 336.555 0.46 ;
    RECT 333.75 0.0 334.375 0.46 ;
    RECT 332.46 0.0 333.47 0.46 ;
    RECT 331.6 0.0 332.18 0.46 ;
    RECT 328.48 0.0 331.32 0.46 ;
    RECT 327.55 0.0 327.85 0.46 ;
    RECT 325.4 0.0 326.975 0.46 ;
    RECT 322.0 0.0 325.12 0.46 ;
    RECT 321.35 0.0 321.72 0.46 ;
    RECT 320.035 0.0 320.77 0.46 ;
    RECT 319.465 0.0 319.755 0.46 ;
    RECT 315.15 0.0 318.92 0.46 ;
    RECT 313.0 0.0 314.87 0.46 ;
    RECT 310.675 0.0 312.72 0.46 ;
    RECT 308.95 0.0 310.395 0.46 ;
    RECT 306.8 0.0 308.67 0.46 ;
    RECT 303.34 0.0 306.52 0.46 ;
    RECT 302.75 0.0 303.06 0.46 ;
    RECT 300.84 0.0 302.47 0.46 ;
    RECT 299.7 0.0 300.32 0.46 ;
    RECT 297.54 0.0 299.42 0.46 ;
    RECT 296.55 0.0 297.26 0.46 ;
    RECT 294.4 0.0 295.97 0.46 ;
    RECT 293.755 0.0 294.12 0.46 ;
    RECT 290.35 0.0 293.475 0.46 ;
    RECT 287.11 0.0 290.07 0.46 ;
    RECT 283.57 0.0 286.83 0.46 ;
    RECT 283.06 0.0 283.29 0.46 ;
    RECT 281.21 0.0 282.78 0.46 ;
    RECT 279.995 0.0 280.63 0.46 ;
    RECT 277.73 0.0 279.715 0.46 ;
    RECT 276.86 0.0 277.45 0.46 ;
    RECT 274.71 0.0 276.34 0.46 ;
    RECT 274.12 0.0 274.43 0.46 ;
    RECT 271.19 0.0 273.84 0.46 ;
    RECT 270.66 0.0 270.91 0.46 ;
    RECT 268.51 0.0 270.38 0.46 ;
    RECT 264.46 0.0 268.23 0.46 ;
    RECT 262.31 0.0 264.18 0.46 ;
    RECT 260.045 0.0 262.03 0.46 ;
    RECT 258.26 0.0 259.765 0.46 ;
    RECT 256.11 0.0 257.98 0.46 ;
    RECT 254.3 0.0 255.83 0.46 ;
    RECT 252.945 0.0 253.5 0.46 ;
    RECT 252.06 0.0 252.665 0.46 ;
    RECT 249.91 0.0 251.78 0.46 ;
    RECT 248.145 0.0 249.63 0.46 ;
    RECT 247.72 0.0 247.865 0.46 ;
    RECT 246.79 0.0 247.44 0.46 ;
    RECT 245.86 0.0 246.51 0.46 ;
    RECT 245.0 0.0 245.58 0.46 ;
    RECT 243.71 0.0 244.72 0.46 ;
    RECT 242.865 0.0 243.43 0.46 ;
    RECT 240.605 0.0 242.585 0.46 ;
    RECT 239.66 0.0 240.0 0.46 ;
    RECT 238.455 0.0 239.38 0.46 ;
    RECT 237.51 0.0 238.175 0.46 ;
    RECT 235.67 0.0 237.23 0.46 ;
    RECT 233.46 0.0 235.39 0.46 ;
    RECT 231.31 0.0 233.18 0.46 ;
    RECT 227.26 0.0 231.03 0.46 ;
    RECT 225.98 0.0 226.98 0.46 ;
    RECT 225.11 0.0 225.7 0.46 ;
    RECT 222.925 0.0 224.83 0.46 ;
    RECT 221.06 0.0 222.645 0.46 ;
    RECT 220.16 0.0 220.52 0.46 ;
    RECT 218.91 0.0 219.88 0.46 ;
    RECT 218.24 0.0 218.63 0.46 ;
    RECT 215.72 0.0 217.96 0.46 ;
    RECT 214.86 0.0 215.44 0.46 ;
    RECT 212.71 0.0 214.58 0.46 ;
    RECT 208.66 0.0 212.43 0.46 ;
    RECT 206.785 0.0 208.38 0.46 ;
    RECT 203.305 0.0 206.23 0.46 ;
    RECT 202.46 0.0 203.025 0.46 ;
    RECT 201.615 0.0 202.18 0.46 ;
    RECT 200.585 0.0 200.995 0.46 ;
    RECT 199.47 0.0 200.03 0.46 ;
    RECT 198.405 0.0 199.19 0.46 ;
    RECT 196.81 0.0 198.125 0.46 ;
    RECT 196.26 0.0 196.53 0.46 ;
    RECT 194.93 0.0 195.72 0.46 ;
    RECT 194.11 0.0 194.65 0.46 ;
    RECT 191.85 0.0 193.83 0.46 ;
    RECT 190.06 0.0 191.57 0.46 ;
    RECT 187.91 0.0 189.78 0.46 ;
    RECT 186.99 0.0 187.63 0.46 ;
    RECT 186.13 0.0 186.71 0.46 ;
    RECT 184.47 0.0 185.85 0.46 ;
    RECT 183.86 0.0 184.19 0.46 ;
    RECT 182.655 0.0 183.295 0.46 ;
    RECT 181.995 0.0 182.375 0.46 ;
    RECT 181.21 0.0 181.43 0.46 ;
    RECT 179.895 0.0 180.565 0.46 ;
    RECT 177.66 0.0 179.265 0.46 ;
    RECT 176.83 0.0 177.085 0.46 ;
    RECT 175.53 0.0 176.55 0.46 ;
    RECT 171.44 0.0 175.25 0.46 ;
    RECT 169.33 0.0 171.16 0.46 ;
    RECT 165.24 0.0 169.05 0.46 ;
    RECT 123.92 0.0 164.96 0.46 ;
    RECT 119.83 0.0 123.64 0.46 ;
    RECT 117.72 0.0 119.55 0.46 ;
    RECT 113.63 0.0 117.44 0.46 ;
    RECT 111.52 0.0 113.35 0.46 ;
    RECT 107.43 0.0 111.24 0.46 ;
    RECT 105.32 0.0 107.15 0.46 ;
    RECT 101.23 0.0 105.04 0.46 ;
    RECT 99.12 0.0 100.95 0.46 ;
    RECT 95.03 0.0 98.84 0.46 ;
    RECT 92.92 0.0 94.75 0.46 ;
    RECT 88.83 0.0 92.64 0.46 ;
    RECT 86.72 0.0 88.55 0.46 ;
    RECT 82.63 0.0 86.44 0.46 ;
    RECT 80.52 0.0 82.35 0.46 ;
    RECT 76.43 0.0 80.24 0.46 ;
    RECT 74.32 0.0 76.15 0.46 ;
    RECT 70.23 0.0 74.04 0.46 ;
    RECT 68.12 0.0 69.95 0.46 ;
    RECT 64.03 0.0 67.84 0.46 ;
    RECT 61.92 0.0 63.75 0.46 ;
    RECT 57.83 0.0 61.64 0.46 ;
    RECT 55.72 0.0 57.55 0.46 ;
    RECT 51.63 0.0 55.44 0.46 ;
    RECT 49.52 0.0 51.35 0.46 ;
    RECT 45.43 0.0 49.24 0.46 ;
    RECT 43.32 0.0 45.15 0.46 ;
    RECT 39.23 0.0 43.04 0.46 ;
    RECT 37.12 0.0 38.95 0.46 ;
    RECT 33.03 0.0 36.84 0.46 ;
    RECT 30.92 0.0 32.75 0.46 ;
    RECT 26.83 0.0 30.64 0.46 ;
    RECT 24.72 0.0 26.55 0.46 ;
    RECT 20.63 0.0 24.44 0.46 ;
    RECT 18.52 0.0 20.35 0.46 ;
    RECT 14.43 0.0 18.24 0.46 ;
    RECT 12.32 0.0 14.15 0.46 ;
    RECT 8.23 0.0 12.04 0.46 ;
    RECT 6.12 0.0 7.95 0.46 ;
    RECT 2.03 0.0 5.84 0.46 ;
    RECT 0.0 0.0 1.75 0.46 ;
    RECT 0.0 0.46 577.18 270.08 ;
    LAYER VIA1 ;
    RECT 0.0 0.0 577.18 270.08 ;
    LAYER M2 DESIGNRULEWIDTH 0.07 ;
    RECT 575.43 0.0 577.18 0.46 ;
    RECT 571.34 0.0 575.15 0.46 ;
    RECT 569.23 0.0 571.06 0.46 ;
    RECT 565.14 0.0 568.95 0.46 ;
    RECT 563.03 0.0 564.86 0.46 ;
    RECT 558.94 0.0 562.75 0.46 ;
    RECT 556.83 0.0 558.66 0.46 ;
    RECT 552.74 0.0 556.55 0.46 ;
    RECT 550.63 0.0 552.46 0.46 ;
    RECT 546.54 0.0 550.35 0.46 ;
    RECT 544.43 0.0 546.26 0.46 ;
    RECT 540.34 0.0 544.15 0.46 ;
    RECT 538.23 0.0 540.06 0.46 ;
    RECT 534.14 0.0 537.95 0.46 ;
    RECT 532.03 0.0 533.86 0.46 ;
    RECT 527.94 0.0 531.75 0.46 ;
    RECT 525.83 0.0 527.66 0.46 ;
    RECT 521.74 0.0 525.55 0.46 ;
    RECT 519.63 0.0 521.46 0.46 ;
    RECT 515.54 0.0 519.35 0.46 ;
    RECT 513.43 0.0 515.26 0.46 ;
    RECT 509.34 0.0 513.15 0.46 ;
    RECT 507.23 0.0 509.06 0.46 ;
    RECT 503.14 0.0 506.95 0.46 ;
    RECT 501.03 0.0 502.86 0.46 ;
    RECT 496.94 0.0 500.75 0.46 ;
    RECT 494.83 0.0 496.66 0.46 ;
    RECT 490.74 0.0 494.55 0.46 ;
    RECT 488.63 0.0 490.46 0.46 ;
    RECT 484.54 0.0 488.35 0.46 ;
    RECT 482.43 0.0 484.26 0.46 ;
    RECT 478.34 0.0 482.15 0.46 ;
    RECT 476.23 0.0 478.06 0.46 ;
    RECT 472.14 0.0 475.95 0.46 ;
    RECT 470.03 0.0 471.86 0.46 ;
    RECT 465.94 0.0 469.75 0.46 ;
    RECT 463.83 0.0 465.66 0.46 ;
    RECT 459.74 0.0 463.55 0.46 ;
    RECT 457.63 0.0 459.46 0.46 ;
    RECT 453.54 0.0 457.35 0.46 ;
    RECT 412.22 0.0 453.26 0.46 ;
    RECT 408.13 0.0 411.94 0.46 ;
    RECT 406.02 0.0 407.85 0.46 ;
    RECT 401.93 0.0 405.74 0.46 ;
    RECT 400.63 0.0 401.65 0.46 ;
    RECT 400.085 0.0 400.35 0.46 ;
    RECT 397.65 0.0 399.52 0.46 ;
    RECT 396.72 0.0 397.37 0.46 ;
    RECT 395.75 0.0 396.17 0.46 ;
    RECT 394.885 0.0 395.17 0.46 ;
    RECT 393.865 0.0 394.265 0.46 ;
    RECT 392.96 0.0 393.32 0.46 ;
    RECT 391.325 0.0 392.68 0.46 ;
    RECT 390.47 0.0 391.045 0.46 ;
    RECT 389.55 0.0 390.19 0.46 ;
    RECT 387.4 0.0 389.27 0.46 ;
    RECT 385.61 0.0 387.12 0.46 ;
    RECT 383.35 0.0 385.33 0.46 ;
    RECT 382.53 0.0 383.07 0.46 ;
    RECT 381.475 0.0 382.25 0.46 ;
    RECT 380.66 0.0 380.92 0.46 ;
    RECT 378.92 0.0 380.38 0.46 ;
    RECT 377.99 0.0 378.64 0.46 ;
    RECT 377.15 0.0 377.71 0.46 ;
    RECT 376.305 0.0 376.87 0.46 ;
    RECT 375.0 0.0 375.505 0.46 ;
    RECT 374.19 0.0 374.72 0.46 ;
    RECT 370.95 0.0 373.91 0.46 ;
    RECT 368.8 0.0 370.385 0.46 ;
    RECT 364.75 0.0 368.52 0.46 ;
    RECT 362.6 0.0 364.47 0.46 ;
    RECT 361.74 0.0 362.32 0.46 ;
    RECT 359.22 0.0 361.46 0.46 ;
    RECT 358.55 0.0 358.94 0.46 ;
    RECT 357.34 0.0 358.27 0.46 ;
    RECT 356.725 0.0 357.06 0.46 ;
    RECT 355.795 0.0 356.12 0.46 ;
    RECT 354.53 0.0 355.515 0.46 ;
    RECT 352.35 0.0 354.25 0.46 ;
    RECT 351.555 0.0 352.07 0.46 ;
    RECT 350.2 0.0 351.275 0.46 ;
    RECT 346.15 0.0 349.92 0.46 ;
    RECT 344.0 0.0 345.87 0.46 ;
    RECT 341.79 0.0 343.72 0.46 ;
    RECT 339.95 0.0 341.51 0.46 ;
    RECT 338.955 0.0 339.67 0.46 ;
    RECT 338.065 0.0 338.675 0.46 ;
    RECT 336.835 0.0 337.52 0.46 ;
    RECT 334.655 0.0 336.555 0.46 ;
    RECT 333.75 0.0 334.375 0.46 ;
    RECT 332.46 0.0 333.47 0.46 ;
    RECT 331.6 0.0 332.18 0.46 ;
    RECT 328.48 0.0 331.32 0.46 ;
    RECT 327.55 0.0 327.85 0.46 ;
    RECT 325.4 0.0 326.975 0.46 ;
    RECT 322.0 0.0 325.12 0.46 ;
    RECT 321.35 0.0 321.72 0.46 ;
    RECT 320.035 0.0 320.77 0.46 ;
    RECT 319.465 0.0 319.755 0.46 ;
    RECT 315.15 0.0 318.92 0.46 ;
    RECT 313.0 0.0 314.87 0.46 ;
    RECT 310.675 0.0 312.72 0.46 ;
    RECT 308.95 0.0 310.395 0.46 ;
    RECT 306.8 0.0 308.67 0.46 ;
    RECT 303.34 0.0 306.52 0.46 ;
    RECT 302.75 0.0 303.06 0.46 ;
    RECT 300.84 0.0 302.47 0.46 ;
    RECT 299.7 0.0 300.32 0.46 ;
    RECT 297.54 0.0 299.42 0.46 ;
    RECT 296.55 0.0 297.26 0.46 ;
    RECT 294.4 0.0 295.97 0.46 ;
    RECT 293.755 0.0 294.12 0.46 ;
    RECT 290.35 0.0 293.475 0.46 ;
    RECT 287.11 0.0 290.07 0.46 ;
    RECT 283.57 0.0 286.83 0.46 ;
    RECT 283.06 0.0 283.29 0.46 ;
    RECT 281.21 0.0 282.78 0.46 ;
    RECT 279.995 0.0 280.63 0.46 ;
    RECT 277.73 0.0 279.715 0.46 ;
    RECT 276.86 0.0 277.45 0.46 ;
    RECT 274.71 0.0 276.34 0.46 ;
    RECT 274.12 0.0 274.43 0.46 ;
    RECT 271.19 0.0 273.84 0.46 ;
    RECT 270.66 0.0 270.91 0.46 ;
    RECT 268.51 0.0 270.38 0.46 ;
    RECT 264.46 0.0 268.23 0.46 ;
    RECT 262.31 0.0 264.18 0.46 ;
    RECT 260.045 0.0 262.03 0.46 ;
    RECT 258.26 0.0 259.765 0.46 ;
    RECT 256.11 0.0 257.98 0.46 ;
    RECT 254.3 0.0 255.83 0.46 ;
    RECT 252.945 0.0 253.5 0.46 ;
    RECT 252.06 0.0 252.665 0.46 ;
    RECT 249.91 0.0 251.78 0.46 ;
    RECT 248.145 0.0 249.63 0.46 ;
    RECT 247.72 0.0 247.865 0.46 ;
    RECT 246.79 0.0 247.44 0.46 ;
    RECT 245.86 0.0 246.51 0.46 ;
    RECT 245.0 0.0 245.58 0.46 ;
    RECT 243.71 0.0 244.72 0.46 ;
    RECT 242.865 0.0 243.43 0.46 ;
    RECT 240.605 0.0 242.585 0.46 ;
    RECT 239.66 0.0 240.0 0.46 ;
    RECT 238.455 0.0 239.38 0.46 ;
    RECT 237.51 0.0 238.175 0.46 ;
    RECT 235.67 0.0 237.23 0.46 ;
    RECT 233.46 0.0 235.39 0.46 ;
    RECT 231.31 0.0 233.18 0.46 ;
    RECT 227.26 0.0 231.03 0.46 ;
    RECT 225.98 0.0 226.98 0.46 ;
    RECT 225.11 0.0 225.7 0.46 ;
    RECT 222.925 0.0 224.83 0.46 ;
    RECT 221.06 0.0 222.645 0.46 ;
    RECT 220.16 0.0 220.52 0.46 ;
    RECT 218.91 0.0 219.88 0.46 ;
    RECT 218.24 0.0 218.63 0.46 ;
    RECT 215.72 0.0 217.96 0.46 ;
    RECT 214.86 0.0 215.44 0.46 ;
    RECT 212.71 0.0 214.58 0.46 ;
    RECT 208.66 0.0 212.43 0.46 ;
    RECT 206.785 0.0 208.38 0.46 ;
    RECT 203.305 0.0 206.23 0.46 ;
    RECT 202.46 0.0 203.025 0.46 ;
    RECT 201.615 0.0 202.18 0.46 ;
    RECT 200.585 0.0 200.995 0.46 ;
    RECT 199.47 0.0 200.03 0.46 ;
    RECT 198.405 0.0 199.19 0.46 ;
    RECT 196.81 0.0 198.125 0.46 ;
    RECT 196.26 0.0 196.53 0.46 ;
    RECT 194.93 0.0 195.72 0.46 ;
    RECT 194.11 0.0 194.65 0.46 ;
    RECT 191.85 0.0 193.83 0.46 ;
    RECT 190.06 0.0 191.57 0.46 ;
    RECT 187.91 0.0 189.78 0.46 ;
    RECT 186.99 0.0 187.63 0.46 ;
    RECT 186.13 0.0 186.71 0.46 ;
    RECT 184.47 0.0 185.85 0.46 ;
    RECT 183.86 0.0 184.19 0.46 ;
    RECT 182.655 0.0 183.295 0.46 ;
    RECT 181.995 0.0 182.375 0.46 ;
    RECT 181.21 0.0 181.43 0.46 ;
    RECT 179.895 0.0 180.565 0.46 ;
    RECT 177.66 0.0 179.265 0.46 ;
    RECT 176.83 0.0 177.085 0.46 ;
    RECT 175.53 0.0 176.55 0.46 ;
    RECT 171.44 0.0 175.25 0.46 ;
    RECT 169.33 0.0 171.16 0.46 ;
    RECT 165.24 0.0 169.05 0.46 ;
    RECT 123.92 0.0 164.96 0.46 ;
    RECT 119.83 0.0 123.64 0.46 ;
    RECT 117.72 0.0 119.55 0.46 ;
    RECT 113.63 0.0 117.44 0.46 ;
    RECT 111.52 0.0 113.35 0.46 ;
    RECT 107.43 0.0 111.24 0.46 ;
    RECT 105.32 0.0 107.15 0.46 ;
    RECT 101.23 0.0 105.04 0.46 ;
    RECT 99.12 0.0 100.95 0.46 ;
    RECT 95.03 0.0 98.84 0.46 ;
    RECT 92.92 0.0 94.75 0.46 ;
    RECT 88.83 0.0 92.64 0.46 ;
    RECT 86.72 0.0 88.55 0.46 ;
    RECT 82.63 0.0 86.44 0.46 ;
    RECT 80.52 0.0 82.35 0.46 ;
    RECT 76.43 0.0 80.24 0.46 ;
    RECT 74.32 0.0 76.15 0.46 ;
    RECT 70.23 0.0 74.04 0.46 ;
    RECT 68.12 0.0 69.95 0.46 ;
    RECT 64.03 0.0 67.84 0.46 ;
    RECT 61.92 0.0 63.75 0.46 ;
    RECT 57.83 0.0 61.64 0.46 ;
    RECT 55.72 0.0 57.55 0.46 ;
    RECT 51.63 0.0 55.44 0.46 ;
    RECT 49.52 0.0 51.35 0.46 ;
    RECT 45.43 0.0 49.24 0.46 ;
    RECT 43.32 0.0 45.15 0.46 ;
    RECT 39.23 0.0 43.04 0.46 ;
    RECT 37.12 0.0 38.95 0.46 ;
    RECT 33.03 0.0 36.84 0.46 ;
    RECT 30.92 0.0 32.75 0.46 ;
    RECT 26.83 0.0 30.64 0.46 ;
    RECT 24.72 0.0 26.55 0.46 ;
    RECT 20.63 0.0 24.44 0.46 ;
    RECT 18.52 0.0 20.35 0.46 ;
    RECT 14.43 0.0 18.24 0.46 ;
    RECT 12.32 0.0 14.15 0.46 ;
    RECT 8.23 0.0 12.04 0.46 ;
    RECT 6.12 0.0 7.95 0.46 ;
    RECT 2.03 0.0 5.84 0.46 ;
    RECT 0.0 0.0 1.75 0.46 ;
    RECT 0.0 0.46 577.18 270.08 ;
    LAYER VIA2 ;
    RECT 0.0 0.0 577.18 270.08 ;
    LAYER M3 DESIGNRULEWIDTH 0.07 ;
    RECT 576.21 0.0 577.18 0.46 ;
    RECT 574.66 0.0 575.645 0.46 ;
    RECT 573.67 0.0 574.38 0.46 ;
    RECT 573.1 0.0 573.39 0.46 ;
    RECT 572.11 0.0 572.82 0.46 ;
    RECT 570.85 0.0 571.83 0.46 ;
    RECT 570.01 0.0 570.32 0.46 ;
    RECT 568.46 0.0 569.445 0.46 ;
    RECT 567.47 0.0 568.18 0.46 ;
    RECT 566.9 0.0 567.19 0.46 ;
    RECT 565.91 0.0 566.62 0.46 ;
    RECT 564.65 0.0 565.63 0.46 ;
    RECT 563.81 0.0 564.12 0.46 ;
    RECT 562.26 0.0 563.245 0.46 ;
    RECT 561.27 0.0 561.98 0.46 ;
    RECT 560.7 0.0 560.99 0.46 ;
    RECT 559.71 0.0 560.42 0.46 ;
    RECT 558.45 0.0 559.43 0.46 ;
    RECT 557.61 0.0 557.92 0.46 ;
    RECT 556.06 0.0 557.045 0.46 ;
    RECT 555.07 0.0 555.78 0.46 ;
    RECT 554.5 0.0 554.79 0.46 ;
    RECT 553.51 0.0 554.22 0.46 ;
    RECT 552.25 0.0 553.23 0.46 ;
    RECT 551.41 0.0 551.72 0.46 ;
    RECT 549.86 0.0 550.845 0.46 ;
    RECT 548.87 0.0 549.58 0.46 ;
    RECT 548.3 0.0 548.59 0.46 ;
    RECT 547.31 0.0 548.02 0.46 ;
    RECT 546.05 0.0 547.03 0.46 ;
    RECT 545.21 0.0 545.52 0.46 ;
    RECT 543.66 0.0 544.645 0.46 ;
    RECT 542.67 0.0 543.38 0.46 ;
    RECT 542.1 0.0 542.39 0.46 ;
    RECT 541.11 0.0 541.82 0.46 ;
    RECT 539.85 0.0 540.83 0.46 ;
    RECT 539.01 0.0 539.32 0.46 ;
    RECT 537.46 0.0 538.445 0.46 ;
    RECT 536.47 0.0 537.18 0.46 ;
    RECT 535.9 0.0 536.19 0.46 ;
    RECT 534.91 0.0 535.62 0.46 ;
    RECT 533.65 0.0 534.63 0.46 ;
    RECT 532.81 0.0 533.12 0.46 ;
    RECT 531.26 0.0 532.245 0.46 ;
    RECT 530.27 0.0 530.98 0.46 ;
    RECT 529.7 0.0 529.99 0.46 ;
    RECT 528.71 0.0 529.42 0.46 ;
    RECT 527.45 0.0 528.43 0.46 ;
    RECT 526.61 0.0 526.92 0.46 ;
    RECT 525.06 0.0 526.045 0.46 ;
    RECT 524.07 0.0 524.78 0.46 ;
    RECT 523.5 0.0 523.79 0.46 ;
    RECT 522.51 0.0 523.22 0.46 ;
    RECT 521.25 0.0 522.23 0.46 ;
    RECT 520.41 0.0 520.72 0.46 ;
    RECT 518.86 0.0 519.845 0.46 ;
    RECT 517.87 0.0 518.58 0.46 ;
    RECT 517.3 0.0 517.59 0.46 ;
    RECT 516.31 0.0 517.02 0.46 ;
    RECT 515.05 0.0 516.03 0.46 ;
    RECT 514.21 0.0 514.52 0.46 ;
    RECT 512.66 0.0 513.645 0.46 ;
    RECT 511.67 0.0 512.38 0.46 ;
    RECT 511.1 0.0 511.39 0.46 ;
    RECT 510.11 0.0 510.82 0.46 ;
    RECT 508.85 0.0 509.83 0.46 ;
    RECT 508.01 0.0 508.32 0.46 ;
    RECT 506.46 0.0 507.445 0.46 ;
    RECT 505.47 0.0 506.18 0.46 ;
    RECT 504.9 0.0 505.19 0.46 ;
    RECT 503.91 0.0 504.62 0.46 ;
    RECT 502.65 0.0 503.63 0.46 ;
    RECT 501.81 0.0 502.12 0.46 ;
    RECT 500.26 0.0 501.245 0.46 ;
    RECT 499.27 0.0 499.98 0.46 ;
    RECT 498.7 0.0 498.99 0.46 ;
    RECT 497.71 0.0 498.42 0.46 ;
    RECT 496.45 0.0 497.43 0.46 ;
    RECT 495.61 0.0 495.92 0.46 ;
    RECT 494.06 0.0 495.045 0.46 ;
    RECT 493.07 0.0 493.78 0.46 ;
    RECT 492.5 0.0 492.79 0.46 ;
    RECT 491.51 0.0 492.22 0.46 ;
    RECT 490.25 0.0 491.23 0.46 ;
    RECT 489.41 0.0 489.72 0.46 ;
    RECT 487.86 0.0 488.845 0.46 ;
    RECT 486.87 0.0 487.58 0.46 ;
    RECT 486.3 0.0 486.59 0.46 ;
    RECT 485.31 0.0 486.02 0.46 ;
    RECT 484.05 0.0 485.03 0.46 ;
    RECT 483.21 0.0 483.52 0.46 ;
    RECT 481.66 0.0 482.645 0.46 ;
    RECT 480.67 0.0 481.38 0.46 ;
    RECT 480.1 0.0 480.39 0.46 ;
    RECT 479.11 0.0 479.82 0.46 ;
    RECT 477.85 0.0 478.83 0.46 ;
    RECT 477.01 0.0 477.32 0.46 ;
    RECT 475.46 0.0 476.445 0.46 ;
    RECT 474.47 0.0 475.18 0.46 ;
    RECT 473.9 0.0 474.19 0.46 ;
    RECT 472.91 0.0 473.62 0.46 ;
    RECT 471.65 0.0 472.63 0.46 ;
    RECT 470.81 0.0 471.12 0.46 ;
    RECT 469.26 0.0 470.245 0.46 ;
    RECT 468.27 0.0 468.98 0.46 ;
    RECT 467.7 0.0 467.99 0.46 ;
    RECT 466.71 0.0 467.42 0.46 ;
    RECT 465.45 0.0 466.43 0.46 ;
    RECT 464.61 0.0 464.92 0.46 ;
    RECT 463.06 0.0 464.045 0.46 ;
    RECT 462.07 0.0 462.78 0.46 ;
    RECT 461.5 0.0 461.79 0.46 ;
    RECT 460.51 0.0 461.22 0.46 ;
    RECT 459.25 0.0 460.23 0.46 ;
    RECT 458.41 0.0 458.72 0.46 ;
    RECT 456.86 0.0 457.845 0.46 ;
    RECT 455.87 0.0 456.58 0.46 ;
    RECT 455.3 0.0 455.59 0.46 ;
    RECT 454.31 0.0 455.02 0.46 ;
    RECT 453.05 0.0 454.03 0.46 ;
    RECT 413.0 0.0 452.52 0.46 ;
    RECT 411.45 0.0 412.435 0.46 ;
    RECT 410.46 0.0 411.17 0.46 ;
    RECT 409.89 0.0 410.18 0.46 ;
    RECT 408.9 0.0 409.61 0.46 ;
    RECT 407.64 0.0 408.62 0.46 ;
    RECT 406.8 0.0 407.11 0.46 ;
    RECT 405.25 0.0 406.235 0.46 ;
    RECT 404.26 0.0 404.97 0.46 ;
    RECT 403.69 0.0 403.98 0.46 ;
    RECT 402.7 0.0 403.41 0.46 ;
    RECT 401.44 0.0 402.42 0.46 ;
    RECT 400.59 0.0 400.91 0.46 ;
    RECT 399.05 0.0 400.07 0.46 ;
    RECT 398.06 0.0 398.77 0.46 ;
    RECT 397.49 0.0 397.78 0.46 ;
    RECT 396.5 0.0 397.21 0.46 ;
    RECT 395.2 0.0 396.22 0.46 ;
    RECT 394.39 0.0 394.68 0.46 ;
    RECT 392.85 0.0 393.87 0.46 ;
    RECT 391.86 0.0 392.57 0.46 ;
    RECT 391.29 0.0 391.58 0.46 ;
    RECT 390.3 0.0 391.01 0.46 ;
    RECT 389.0 0.0 390.02 0.46 ;
    RECT 388.19 0.0 388.48 0.46 ;
    RECT 386.65 0.0 387.67 0.46 ;
    RECT 385.66 0.0 386.37 0.46 ;
    RECT 385.09 0.0 385.38 0.46 ;
    RECT 384.1 0.0 384.81 0.46 ;
    RECT 382.8 0.0 383.82 0.46 ;
    RECT 381.99 0.0 382.28 0.46 ;
    RECT 380.45 0.0 381.47 0.46 ;
    RECT 379.46 0.0 380.17 0.46 ;
    RECT 378.89 0.0 379.18 0.46 ;
    RECT 377.9 0.0 378.61 0.46 ;
    RECT 376.6 0.0 377.62 0.46 ;
    RECT 375.79 0.0 376.08 0.46 ;
    RECT 374.25 0.0 375.27 0.46 ;
    RECT 373.26 0.0 373.97 0.46 ;
    RECT 372.69 0.0 372.98 0.46 ;
    RECT 371.7 0.0 372.41 0.46 ;
    RECT 370.4 0.0 371.42 0.46 ;
    RECT 369.59 0.0 369.88 0.46 ;
    RECT 368.05 0.0 369.07 0.46 ;
    RECT 367.06 0.0 367.77 0.46 ;
    RECT 366.49 0.0 366.78 0.46 ;
    RECT 365.5 0.0 366.21 0.46 ;
    RECT 364.2 0.0 365.22 0.46 ;
    RECT 363.39 0.0 363.68 0.46 ;
    RECT 361.85 0.0 362.87 0.46 ;
    RECT 360.86 0.0 361.57 0.46 ;
    RECT 360.29 0.0 360.58 0.46 ;
    RECT 359.3 0.0 360.01 0.46 ;
    RECT 358.0 0.0 359.02 0.46 ;
    RECT 357.19 0.0 357.48 0.46 ;
    RECT 355.65 0.0 356.67 0.46 ;
    RECT 354.66 0.0 355.37 0.46 ;
    RECT 354.09 0.0 354.38 0.46 ;
    RECT 353.1 0.0 353.81 0.46 ;
    RECT 351.8 0.0 352.82 0.46 ;
    RECT 350.99 0.0 351.28 0.46 ;
    RECT 349.45 0.0 350.47 0.46 ;
    RECT 348.46 0.0 349.17 0.46 ;
    RECT 347.89 0.0 348.18 0.46 ;
    RECT 346.9 0.0 347.61 0.46 ;
    RECT 345.6 0.0 346.62 0.46 ;
    RECT 344.79 0.0 345.08 0.46 ;
    RECT 343.25 0.0 344.27 0.46 ;
    RECT 342.26 0.0 342.97 0.46 ;
    RECT 341.69 0.0 341.98 0.46 ;
    RECT 340.7 0.0 341.41 0.46 ;
    RECT 339.4 0.0 340.42 0.46 ;
    RECT 338.59 0.0 338.88 0.46 ;
    RECT 337.05 0.0 338.07 0.46 ;
    RECT 336.06 0.0 336.77 0.46 ;
    RECT 335.49 0.0 335.78 0.46 ;
    RECT 334.5 0.0 335.21 0.46 ;
    RECT 333.2 0.0 334.22 0.46 ;
    RECT 332.39 0.0 332.68 0.46 ;
    RECT 330.85 0.0 331.87 0.46 ;
    RECT 329.86 0.0 330.57 0.46 ;
    RECT 329.29 0.0 329.58 0.46 ;
    RECT 328.3 0.0 329.01 0.46 ;
    RECT 327.0 0.0 328.02 0.46 ;
    RECT 326.19 0.0 326.48 0.46 ;
    RECT 324.65 0.0 325.67 0.46 ;
    RECT 323.66 0.0 324.37 0.46 ;
    RECT 323.09 0.0 323.38 0.46 ;
    RECT 322.1 0.0 322.81 0.46 ;
    RECT 320.8 0.0 321.82 0.46 ;
    RECT 319.99 0.0 320.28 0.46 ;
    RECT 318.45 0.0 319.47 0.46 ;
    RECT 317.46 0.0 318.17 0.46 ;
    RECT 316.89 0.0 317.18 0.46 ;
    RECT 315.9 0.0 316.61 0.46 ;
    RECT 314.6 0.0 315.62 0.46 ;
    RECT 313.79 0.0 314.08 0.46 ;
    RECT 312.25 0.0 313.27 0.46 ;
    RECT 311.26 0.0 311.97 0.46 ;
    RECT 310.69 0.0 310.98 0.46 ;
    RECT 309.7 0.0 310.41 0.46 ;
    RECT 308.4 0.0 309.42 0.46 ;
    RECT 307.59 0.0 307.88 0.46 ;
    RECT 306.05 0.0 307.07 0.46 ;
    RECT 305.06 0.0 305.77 0.46 ;
    RECT 304.49 0.0 304.78 0.46 ;
    RECT 303.5 0.0 304.21 0.46 ;
    RECT 302.2 0.0 303.22 0.46 ;
    RECT 301.39 0.0 301.68 0.46 ;
    RECT 299.85 0.0 300.87 0.46 ;
    RECT 298.86 0.0 299.57 0.46 ;
    RECT 298.29 0.0 298.58 0.46 ;
    RECT 297.3 0.0 298.01 0.46 ;
    RECT 296.0 0.0 297.02 0.46 ;
    RECT 295.19 0.0 295.48 0.46 ;
    RECT 293.65 0.0 294.67 0.46 ;
    RECT 292.66 0.0 293.37 0.46 ;
    RECT 292.09 0.0 292.38 0.46 ;
    RECT 291.1 0.0 291.81 0.46 ;
    RECT 289.8 0.0 290.82 0.46 ;
    RECT 287.9 0.0 289.28 0.46 ;
    RECT 286.36 0.0 287.38 0.46 ;
    RECT 285.37 0.0 286.08 0.46 ;
    RECT 284.8 0.0 285.09 0.46 ;
    RECT 283.81 0.0 284.52 0.46 ;
    RECT 282.51 0.0 283.53 0.46 ;
    RECT 281.7 0.0 281.99 0.46 ;
    RECT 280.16 0.0 281.18 0.46 ;
    RECT 279.17 0.0 279.88 0.46 ;
    RECT 278.6 0.0 278.89 0.46 ;
    RECT 277.61 0.0 278.32 0.46 ;
    RECT 276.31 0.0 277.33 0.46 ;
    RECT 275.5 0.0 275.79 0.46 ;
    RECT 273.96 0.0 274.98 0.46 ;
    RECT 272.97 0.0 273.68 0.46 ;
    RECT 272.4 0.0 272.69 0.46 ;
    RECT 271.41 0.0 272.12 0.46 ;
    RECT 270.11 0.0 271.13 0.46 ;
    RECT 269.3 0.0 269.59 0.46 ;
    RECT 267.76 0.0 268.78 0.46 ;
    RECT 266.77 0.0 267.48 0.46 ;
    RECT 266.2 0.0 266.49 0.46 ;
    RECT 265.21 0.0 265.92 0.46 ;
    RECT 263.91 0.0 264.93 0.46 ;
    RECT 263.1 0.0 263.39 0.46 ;
    RECT 261.56 0.0 262.58 0.46 ;
    RECT 260.57 0.0 261.28 0.46 ;
    RECT 260.0 0.0 260.29 0.46 ;
    RECT 259.01 0.0 259.72 0.46 ;
    RECT 257.71 0.0 258.73 0.46 ;
    RECT 256.9 0.0 257.19 0.46 ;
    RECT 255.36 0.0 256.38 0.46 ;
    RECT 254.37 0.0 255.08 0.46 ;
    RECT 253.8 0.0 254.09 0.46 ;
    RECT 252.81 0.0 253.52 0.46 ;
    RECT 251.51 0.0 252.53 0.46 ;
    RECT 250.7 0.0 250.99 0.46 ;
    RECT 249.16 0.0 250.18 0.46 ;
    RECT 248.17 0.0 248.88 0.46 ;
    RECT 247.6 0.0 247.89 0.46 ;
    RECT 246.61 0.0 247.32 0.46 ;
    RECT 245.31 0.0 246.33 0.46 ;
    RECT 244.5 0.0 244.79 0.46 ;
    RECT 242.96 0.0 243.98 0.46 ;
    RECT 241.97 0.0 242.68 0.46 ;
    RECT 241.4 0.0 241.69 0.46 ;
    RECT 240.41 0.0 241.12 0.46 ;
    RECT 239.11 0.0 240.13 0.46 ;
    RECT 238.3 0.0 238.59 0.46 ;
    RECT 236.76 0.0 237.78 0.46 ;
    RECT 235.77 0.0 236.48 0.46 ;
    RECT 235.2 0.0 235.49 0.46 ;
    RECT 234.21 0.0 234.92 0.46 ;
    RECT 232.91 0.0 233.93 0.46 ;
    RECT 232.1 0.0 232.39 0.46 ;
    RECT 230.56 0.0 231.58 0.46 ;
    RECT 229.57 0.0 230.28 0.46 ;
    RECT 229.0 0.0 229.29 0.46 ;
    RECT 228.01 0.0 228.72 0.46 ;
    RECT 226.71 0.0 227.73 0.46 ;
    RECT 225.9 0.0 226.19 0.46 ;
    RECT 224.36 0.0 225.38 0.46 ;
    RECT 223.37 0.0 224.08 0.46 ;
    RECT 222.8 0.0 223.09 0.46 ;
    RECT 221.81 0.0 222.52 0.46 ;
    RECT 220.51 0.0 221.53 0.46 ;
    RECT 219.7 0.0 219.99 0.46 ;
    RECT 218.16 0.0 219.18 0.46 ;
    RECT 217.17 0.0 217.88 0.46 ;
    RECT 216.6 0.0 216.89 0.46 ;
    RECT 215.61 0.0 216.32 0.46 ;
    RECT 214.31 0.0 215.33 0.46 ;
    RECT 213.5 0.0 213.79 0.46 ;
    RECT 211.96 0.0 212.98 0.46 ;
    RECT 210.97 0.0 211.68 0.46 ;
    RECT 210.4 0.0 210.69 0.46 ;
    RECT 208.11 0.0 210.12 0.46 ;
    RECT 207.3 0.0 207.59 0.46 ;
    RECT 205.76 0.0 206.78 0.46 ;
    RECT 204.77 0.0 205.48 0.46 ;
    RECT 204.2 0.0 204.49 0.46 ;
    RECT 203.21 0.0 203.92 0.46 ;
    RECT 201.91 0.0 202.93 0.46 ;
    RECT 201.1 0.0 201.39 0.46 ;
    RECT 199.56 0.0 200.58 0.46 ;
    RECT 198.57 0.0 199.28 0.46 ;
    RECT 198.0 0.0 198.29 0.46 ;
    RECT 197.01 0.0 197.72 0.46 ;
    RECT 195.71 0.0 196.73 0.46 ;
    RECT 194.9 0.0 195.19 0.46 ;
    RECT 193.36 0.0 194.38 0.46 ;
    RECT 192.37 0.0 193.08 0.46 ;
    RECT 191.8 0.0 192.09 0.46 ;
    RECT 190.81 0.0 191.52 0.46 ;
    RECT 189.51 0.0 190.53 0.46 ;
    RECT 188.7 0.0 188.99 0.46 ;
    RECT 187.16 0.0 188.18 0.46 ;
    RECT 186.17 0.0 186.88 0.46 ;
    RECT 185.6 0.0 185.89 0.46 ;
    RECT 184.61 0.0 185.32 0.46 ;
    RECT 183.31 0.0 184.33 0.46 ;
    RECT 182.5 0.0 182.79 0.46 ;
    RECT 180.96 0.0 181.98 0.46 ;
    RECT 179.97 0.0 180.68 0.46 ;
    RECT 179.4 0.0 179.69 0.46 ;
    RECT 178.41 0.0 179.12 0.46 ;
    RECT 177.11 0.0 178.13 0.46 ;
    RECT 176.27 0.0 176.59 0.46 ;
    RECT 174.76 0.0 175.74 0.46 ;
    RECT 173.77 0.0 174.48 0.46 ;
    RECT 173.2 0.0 173.49 0.46 ;
    RECT 172.21 0.0 172.92 0.46 ;
    RECT 170.945 0.0 171.93 0.46 ;
    RECT 170.07 0.0 170.38 0.46 ;
    RECT 168.56 0.0 169.54 0.46 ;
    RECT 167.57 0.0 168.28 0.46 ;
    RECT 167.0 0.0 167.29 0.46 ;
    RECT 166.01 0.0 166.72 0.46 ;
    RECT 164.745 0.0 165.73 0.46 ;
    RECT 124.66 0.0 164.18 0.46 ;
    RECT 123.15 0.0 124.13 0.46 ;
    RECT 122.16 0.0 122.87 0.46 ;
    RECT 121.59 0.0 121.88 0.46 ;
    RECT 120.6 0.0 121.31 0.46 ;
    RECT 119.335 0.0 120.32 0.46 ;
    RECT 118.46 0.0 118.77 0.46 ;
    RECT 116.95 0.0 117.93 0.46 ;
    RECT 115.96 0.0 116.67 0.46 ;
    RECT 115.39 0.0 115.68 0.46 ;
    RECT 114.4 0.0 115.11 0.46 ;
    RECT 113.135 0.0 114.12 0.46 ;
    RECT 112.26 0.0 112.57 0.46 ;
    RECT 110.75 0.0 111.73 0.46 ;
    RECT 109.76 0.0 110.47 0.46 ;
    RECT 109.19 0.0 109.48 0.46 ;
    RECT 108.2 0.0 108.91 0.46 ;
    RECT 106.935 0.0 107.92 0.46 ;
    RECT 106.06 0.0 106.37 0.46 ;
    RECT 104.55 0.0 105.53 0.46 ;
    RECT 103.56 0.0 104.27 0.46 ;
    RECT 102.99 0.0 103.28 0.46 ;
    RECT 102.0 0.0 102.71 0.46 ;
    RECT 100.735 0.0 101.72 0.46 ;
    RECT 99.86 0.0 100.17 0.46 ;
    RECT 98.35 0.0 99.33 0.46 ;
    RECT 97.36 0.0 98.07 0.46 ;
    RECT 96.79 0.0 97.08 0.46 ;
    RECT 95.8 0.0 96.51 0.46 ;
    RECT 94.535 0.0 95.52 0.46 ;
    RECT 93.66 0.0 93.97 0.46 ;
    RECT 92.15 0.0 93.13 0.46 ;
    RECT 91.16 0.0 91.87 0.46 ;
    RECT 90.59 0.0 90.88 0.46 ;
    RECT 89.6 0.0 90.31 0.46 ;
    RECT 88.335 0.0 89.32 0.46 ;
    RECT 87.46 0.0 87.77 0.46 ;
    RECT 85.95 0.0 86.93 0.46 ;
    RECT 84.96 0.0 85.67 0.46 ;
    RECT 84.39 0.0 84.68 0.46 ;
    RECT 83.4 0.0 84.11 0.46 ;
    RECT 82.135 0.0 83.12 0.46 ;
    RECT 81.26 0.0 81.57 0.46 ;
    RECT 79.75 0.0 80.73 0.46 ;
    RECT 78.76 0.0 79.47 0.46 ;
    RECT 78.19 0.0 78.48 0.46 ;
    RECT 77.2 0.0 77.91 0.46 ;
    RECT 75.935 0.0 76.92 0.46 ;
    RECT 75.06 0.0 75.37 0.46 ;
    RECT 73.55 0.0 74.53 0.46 ;
    RECT 72.56 0.0 73.27 0.46 ;
    RECT 71.99 0.0 72.28 0.46 ;
    RECT 71.0 0.0 71.71 0.46 ;
    RECT 69.735 0.0 70.72 0.46 ;
    RECT 68.86 0.0 69.17 0.46 ;
    RECT 67.35 0.0 68.33 0.46 ;
    RECT 66.36 0.0 67.07 0.46 ;
    RECT 65.79 0.0 66.08 0.46 ;
    RECT 64.8 0.0 65.51 0.46 ;
    RECT 63.535 0.0 64.52 0.46 ;
    RECT 62.66 0.0 62.97 0.46 ;
    RECT 61.15 0.0 62.13 0.46 ;
    RECT 60.16 0.0 60.87 0.46 ;
    RECT 59.59 0.0 59.88 0.46 ;
    RECT 58.6 0.0 59.31 0.46 ;
    RECT 57.335 0.0 58.32 0.46 ;
    RECT 56.46 0.0 56.77 0.46 ;
    RECT 54.95 0.0 55.93 0.46 ;
    RECT 53.96 0.0 54.67 0.46 ;
    RECT 53.39 0.0 53.68 0.46 ;
    RECT 52.4 0.0 53.11 0.46 ;
    RECT 51.135 0.0 52.12 0.46 ;
    RECT 50.26 0.0 50.57 0.46 ;
    RECT 48.75 0.0 49.73 0.46 ;
    RECT 47.76 0.0 48.47 0.46 ;
    RECT 47.19 0.0 47.48 0.46 ;
    RECT 46.2 0.0 46.91 0.46 ;
    RECT 44.935 0.0 45.92 0.46 ;
    RECT 44.06 0.0 44.37 0.46 ;
    RECT 42.55 0.0 43.53 0.46 ;
    RECT 41.56 0.0 42.27 0.46 ;
    RECT 40.99 0.0 41.28 0.46 ;
    RECT 40.0 0.0 40.71 0.46 ;
    RECT 38.735 0.0 39.72 0.46 ;
    RECT 37.86 0.0 38.17 0.46 ;
    RECT 36.35 0.0 37.33 0.46 ;
    RECT 35.36 0.0 36.07 0.46 ;
    RECT 34.79 0.0 35.08 0.46 ;
    RECT 33.8 0.0 34.51 0.46 ;
    RECT 32.535 0.0 33.52 0.46 ;
    RECT 31.66 0.0 31.97 0.46 ;
    RECT 30.15 0.0 31.13 0.46 ;
    RECT 29.16 0.0 29.87 0.46 ;
    RECT 28.59 0.0 28.88 0.46 ;
    RECT 27.6 0.0 28.31 0.46 ;
    RECT 26.335 0.0 27.32 0.46 ;
    RECT 25.46 0.0 25.77 0.46 ;
    RECT 23.95 0.0 24.93 0.46 ;
    RECT 22.96 0.0 23.67 0.46 ;
    RECT 22.39 0.0 22.68 0.46 ;
    RECT 21.4 0.0 22.11 0.46 ;
    RECT 20.135 0.0 21.12 0.46 ;
    RECT 19.26 0.0 19.57 0.46 ;
    RECT 17.75 0.0 18.73 0.46 ;
    RECT 16.76 0.0 17.47 0.46 ;
    RECT 16.19 0.0 16.48 0.46 ;
    RECT 15.2 0.0 15.91 0.46 ;
    RECT 13.935 0.0 14.92 0.46 ;
    RECT 13.06 0.0 13.37 0.46 ;
    RECT 11.55 0.0 12.53 0.46 ;
    RECT 10.56 0.0 11.27 0.46 ;
    RECT 9.99 0.0 10.28 0.46 ;
    RECT 9.0 0.0 9.71 0.46 ;
    RECT 7.735 0.0 8.72 0.46 ;
    RECT 6.86 0.0 7.17 0.46 ;
    RECT 5.35 0.0 6.33 0.46 ;
    RECT 4.36 0.0 5.07 0.46 ;
    RECT 3.79 0.0 4.08 0.46 ;
    RECT 2.8 0.0 3.51 0.46 ;
    RECT 1.535 0.0 2.52 0.46 ;
    RECT 0.0 0.0 0.97 0.46 ;
    RECT 0.0 0.46 577.18 270.08 ;
    LAYER VIA3 ;
    RECT 0.0 0.0 577.18 270.08 ;
    LAYER M4 DESIGNRULEWIDTH 0.07 ;
    RECT 576.8 0.0 577.18 0.46 ;
    RECT 576.45 0.0 576.59 0.46 ;
    RECT 574.9 0.0 575.4 0.46 ;
    RECT 573.67 0.0 574.38 0.46 ;
    RECT 572.11 0.0 572.82 0.46 ;
    RECT 571.09 0.0 571.59 0.46 ;
    RECT 568.7 0.0 569.2 0.46 ;
    RECT 567.47 0.0 568.18 0.46 ;
    RECT 565.91 0.0 566.62 0.46 ;
    RECT 564.89 0.0 565.39 0.46 ;
    RECT 562.5 0.0 563.0 0.46 ;
    RECT 561.27 0.0 561.98 0.46 ;
    RECT 559.71 0.0 560.42 0.46 ;
    RECT 558.69 0.0 559.19 0.46 ;
    RECT 556.3 0.0 556.8 0.46 ;
    RECT 555.07 0.0 555.78 0.46 ;
    RECT 553.51 0.0 554.22 0.46 ;
    RECT 552.49 0.0 552.99 0.46 ;
    RECT 550.1 0.0 550.6 0.46 ;
    RECT 548.87 0.0 549.58 0.46 ;
    RECT 547.31 0.0 548.02 0.46 ;
    RECT 546.29 0.0 546.79 0.46 ;
    RECT 543.9 0.0 544.4 0.46 ;
    RECT 542.67 0.0 543.38 0.46 ;
    RECT 541.11 0.0 541.82 0.46 ;
    RECT 540.09 0.0 540.59 0.46 ;
    RECT 537.7 0.0 538.2 0.46 ;
    RECT 536.47 0.0 537.18 0.46 ;
    RECT 534.91 0.0 535.62 0.46 ;
    RECT 533.89 0.0 534.39 0.46 ;
    RECT 531.5 0.0 532.0 0.46 ;
    RECT 530.27 0.0 530.98 0.46 ;
    RECT 528.71 0.0 529.42 0.46 ;
    RECT 527.69 0.0 528.19 0.46 ;
    RECT 525.3 0.0 525.8 0.46 ;
    RECT 524.07 0.0 524.78 0.46 ;
    RECT 522.51 0.0 523.22 0.46 ;
    RECT 521.49 0.0 521.99 0.46 ;
    RECT 519.1 0.0 519.6 0.46 ;
    RECT 517.87 0.0 518.58 0.46 ;
    RECT 516.31 0.0 517.02 0.46 ;
    RECT 515.29 0.0 515.79 0.46 ;
    RECT 512.9 0.0 513.4 0.46 ;
    RECT 511.67 0.0 512.38 0.46 ;
    RECT 510.11 0.0 510.82 0.46 ;
    RECT 509.09 0.0 509.59 0.46 ;
    RECT 506.7 0.0 507.2 0.46 ;
    RECT 505.47 0.0 506.18 0.46 ;
    RECT 503.91 0.0 504.62 0.46 ;
    RECT 502.89 0.0 503.39 0.46 ;
    RECT 500.5 0.0 501.0 0.46 ;
    RECT 499.27 0.0 499.98 0.46 ;
    RECT 497.71 0.0 498.42 0.46 ;
    RECT 496.69 0.0 497.19 0.46 ;
    RECT 494.3 0.0 494.8 0.46 ;
    RECT 493.07 0.0 493.78 0.46 ;
    RECT 491.51 0.0 492.22 0.46 ;
    RECT 490.49 0.0 490.99 0.46 ;
    RECT 488.1 0.0 488.6 0.46 ;
    RECT 486.87 0.0 487.58 0.46 ;
    RECT 485.31 0.0 486.02 0.46 ;
    RECT 484.29 0.0 484.79 0.46 ;
    RECT 481.9 0.0 482.4 0.46 ;
    RECT 480.67 0.0 481.38 0.46 ;
    RECT 479.11 0.0 479.82 0.46 ;
    RECT 478.09 0.0 478.59 0.46 ;
    RECT 475.7 0.0 476.2 0.46 ;
    RECT 474.47 0.0 475.18 0.46 ;
    RECT 472.91 0.0 473.62 0.46 ;
    RECT 471.89 0.0 472.39 0.46 ;
    RECT 469.5 0.0 470.0 0.46 ;
    RECT 468.27 0.0 468.98 0.46 ;
    RECT 466.71 0.0 467.42 0.46 ;
    RECT 465.69 0.0 466.19 0.46 ;
    RECT 463.3 0.0 463.8 0.46 ;
    RECT 462.07 0.0 462.78 0.46 ;
    RECT 460.51 0.0 461.22 0.46 ;
    RECT 459.49 0.0 459.99 0.46 ;
    RECT 457.1 0.0 457.6 0.46 ;
    RECT 455.87 0.0 456.58 0.46 ;
    RECT 454.31 0.0 455.02 0.46 ;
    RECT 453.29 0.0 453.79 0.46 ;
    RECT 451.115 0.0 452.24 0.46 ;
    RECT 450.725 0.0 450.905 0.46 ;
    RECT 448.845 0.0 450.515 0.46 ;
    RECT 447.78 0.0 448.635 0.46 ;
    RECT 445.12 0.0 447.57 0.46 ;
    RECT 444.8 0.0 444.91 0.46 ;
    RECT 443.135 0.0 444.59 0.46 ;
    RECT 442.815 0.0 442.925 0.46 ;
    RECT 441.01 0.0 442.605 0.46 ;
    RECT 439.675 0.0 440.52 0.46 ;
    RECT 439.355 0.0 439.465 0.46 ;
    RECT 438.655 0.0 439.145 0.46 ;
    RECT 437.765 0.0 438.445 0.46 ;
    RECT 436.705 0.0 437.555 0.46 ;
    RECT 436.385 0.0 436.495 0.46 ;
    RECT 435.475 0.0 436.175 0.46 ;
    RECT 433.44 0.0 435.265 0.46 ;
    RECT 432.25 0.0 433.23 0.46 ;
    RECT 430.215 0.0 432.04 0.46 ;
    RECT 429.305 0.0 430.005 0.46 ;
    RECT 428.985 0.0 429.095 0.46 ;
    RECT 427.925 0.0 428.775 0.46 ;
    RECT 427.035 0.0 427.715 0.46 ;
    RECT 426.335 0.0 426.825 0.46 ;
    RECT 426.015 0.0 426.125 0.46 ;
    RECT 424.68 0.0 425.805 0.46 ;
    RECT 422.875 0.0 424.47 0.46 ;
    RECT 422.555 0.0 422.665 0.46 ;
    RECT 420.89 0.0 422.345 0.46 ;
    RECT 420.57 0.0 420.68 0.46 ;
    RECT 417.91 0.0 420.36 0.46 ;
    RECT 416.845 0.0 417.7 0.46 ;
    RECT 414.965 0.0 416.635 0.46 ;
    RECT 414.575 0.0 414.755 0.46 ;
    RECT 413.24 0.0 414.365 0.46 ;
    RECT 411.69 0.0 412.19 0.46 ;
    RECT 410.46 0.0 411.17 0.46 ;
    RECT 408.9 0.0 409.61 0.46 ;
    RECT 407.88 0.0 408.38 0.46 ;
    RECT 405.49 0.0 405.99 0.46 ;
    RECT 404.26 0.0 404.97 0.46 ;
    RECT 402.7 0.0 403.41 0.46 ;
    RECT 401.68 0.0 402.18 0.46 ;
    RECT 399.29 0.0 399.79 0.46 ;
    RECT 398.06 0.0 398.77 0.46 ;
    RECT 396.5 0.0 397.21 0.46 ;
    RECT 395.48 0.0 395.98 0.46 ;
    RECT 393.09 0.0 393.59 0.46 ;
    RECT 391.86 0.0 392.57 0.46 ;
    RECT 390.3 0.0 391.01 0.46 ;
    RECT 389.28 0.0 389.78 0.46 ;
    RECT 386.89 0.0 387.39 0.46 ;
    RECT 385.66 0.0 386.37 0.46 ;
    RECT 384.1 0.0 384.81 0.46 ;
    RECT 383.08 0.0 383.58 0.46 ;
    RECT 380.69 0.0 381.19 0.46 ;
    RECT 379.46 0.0 380.17 0.46 ;
    RECT 377.9 0.0 378.61 0.46 ;
    RECT 376.88 0.0 377.38 0.46 ;
    RECT 374.49 0.0 374.99 0.46 ;
    RECT 373.26 0.0 373.97 0.46 ;
    RECT 371.7 0.0 372.41 0.46 ;
    RECT 370.68 0.0 371.18 0.46 ;
    RECT 368.29 0.0 368.79 0.46 ;
    RECT 367.06 0.0 367.77 0.46 ;
    RECT 365.5 0.0 366.21 0.46 ;
    RECT 364.48 0.0 364.98 0.46 ;
    RECT 362.09 0.0 362.59 0.46 ;
    RECT 360.86 0.0 361.57 0.46 ;
    RECT 359.3 0.0 360.01 0.46 ;
    RECT 358.28 0.0 358.78 0.46 ;
    RECT 355.89 0.0 356.39 0.46 ;
    RECT 354.66 0.0 355.37 0.46 ;
    RECT 353.1 0.0 353.81 0.46 ;
    RECT 352.08 0.0 352.58 0.46 ;
    RECT 349.69 0.0 350.19 0.46 ;
    RECT 348.46 0.0 349.17 0.46 ;
    RECT 346.9 0.0 347.61 0.46 ;
    RECT 345.88 0.0 346.38 0.46 ;
    RECT 343.49 0.0 343.99 0.46 ;
    RECT 342.26 0.0 342.97 0.46 ;
    RECT 340.7 0.0 341.41 0.46 ;
    RECT 339.68 0.0 340.18 0.46 ;
    RECT 337.29 0.0 337.79 0.46 ;
    RECT 336.06 0.0 336.77 0.46 ;
    RECT 334.5 0.0 335.21 0.46 ;
    RECT 333.48 0.0 333.98 0.46 ;
    RECT 331.09 0.0 331.59 0.46 ;
    RECT 329.86 0.0 330.57 0.46 ;
    RECT 328.3 0.0 329.01 0.46 ;
    RECT 327.28 0.0 327.78 0.46 ;
    RECT 324.89 0.0 325.39 0.46 ;
    RECT 323.66 0.0 324.37 0.46 ;
    RECT 322.1 0.0 322.81 0.46 ;
    RECT 321.08 0.0 321.58 0.46 ;
    RECT 318.69 0.0 319.19 0.46 ;
    RECT 317.46 0.0 318.17 0.46 ;
    RECT 315.9 0.0 316.61 0.46 ;
    RECT 314.88 0.0 315.38 0.46 ;
    RECT 312.49 0.0 312.99 0.46 ;
    RECT 311.26 0.0 311.97 0.46 ;
    RECT 309.7 0.0 310.41 0.46 ;
    RECT 308.68 0.0 309.18 0.46 ;
    RECT 306.29 0.0 306.79 0.46 ;
    RECT 305.06 0.0 305.77 0.46 ;
    RECT 303.5 0.0 304.21 0.46 ;
    RECT 302.48 0.0 302.98 0.46 ;
    RECT 300.09 0.0 300.59 0.46 ;
    RECT 298.86 0.0 299.57 0.46 ;
    RECT 297.3 0.0 298.01 0.46 ;
    RECT 296.28 0.0 296.78 0.46 ;
    RECT 293.89 0.0 294.39 0.46 ;
    RECT 292.66 0.0 293.37 0.46 ;
    RECT 291.1 0.0 291.81 0.46 ;
    RECT 290.08 0.0 290.58 0.46 ;
    RECT 288.15 0.0 289.03 0.46 ;
    RECT 286.6 0.0 287.1 0.46 ;
    RECT 285.37 0.0 286.08 0.46 ;
    RECT 283.81 0.0 284.52 0.46 ;
    RECT 282.79 0.0 283.29 0.46 ;
    RECT 280.4 0.0 280.9 0.46 ;
    RECT 279.17 0.0 279.88 0.46 ;
    RECT 277.61 0.0 278.32 0.46 ;
    RECT 276.59 0.0 277.09 0.46 ;
    RECT 274.2 0.0 274.7 0.46 ;
    RECT 272.97 0.0 273.68 0.46 ;
    RECT 271.41 0.0 272.12 0.46 ;
    RECT 270.39 0.0 270.89 0.46 ;
    RECT 268.0 0.0 268.5 0.46 ;
    RECT 266.77 0.0 267.48 0.46 ;
    RECT 265.21 0.0 265.92 0.46 ;
    RECT 264.19 0.0 264.69 0.46 ;
    RECT 261.8 0.0 262.3 0.46 ;
    RECT 260.57 0.0 261.28 0.46 ;
    RECT 259.01 0.0 259.72 0.46 ;
    RECT 257.99 0.0 258.49 0.46 ;
    RECT 255.6 0.0 256.1 0.46 ;
    RECT 254.37 0.0 255.08 0.46 ;
    RECT 252.81 0.0 253.52 0.46 ;
    RECT 251.79 0.0 252.29 0.46 ;
    RECT 249.4 0.0 249.9 0.46 ;
    RECT 248.17 0.0 248.88 0.46 ;
    RECT 246.61 0.0 247.32 0.46 ;
    RECT 245.59 0.0 246.09 0.46 ;
    RECT 243.2 0.0 243.7 0.46 ;
    RECT 241.97 0.0 242.68 0.46 ;
    RECT 240.41 0.0 241.12 0.46 ;
    RECT 239.39 0.0 239.89 0.46 ;
    RECT 237.0 0.0 237.5 0.46 ;
    RECT 235.77 0.0 236.48 0.46 ;
    RECT 234.21 0.0 234.92 0.46 ;
    RECT 233.19 0.0 233.69 0.46 ;
    RECT 230.8 0.0 231.3 0.46 ;
    RECT 229.57 0.0 230.28 0.46 ;
    RECT 228.01 0.0 228.72 0.46 ;
    RECT 226.99 0.0 227.49 0.46 ;
    RECT 224.6 0.0 225.1 0.46 ;
    RECT 223.37 0.0 224.08 0.46 ;
    RECT 221.81 0.0 222.52 0.46 ;
    RECT 220.79 0.0 221.29 0.46 ;
    RECT 218.4 0.0 218.9 0.46 ;
    RECT 217.17 0.0 217.88 0.46 ;
    RECT 215.61 0.0 216.32 0.46 ;
    RECT 214.59 0.0 215.09 0.46 ;
    RECT 212.2 0.0 212.7 0.46 ;
    RECT 210.97 0.0 211.68 0.46 ;
    RECT 209.41 0.0 210.12 0.46 ;
    RECT 208.39 0.0 208.89 0.46 ;
    RECT 206.0 0.0 206.5 0.46 ;
    RECT 204.77 0.0 205.48 0.46 ;
    RECT 203.21 0.0 203.92 0.46 ;
    RECT 202.19 0.0 202.69 0.46 ;
    RECT 199.8 0.0 200.3 0.46 ;
    RECT 198.57 0.0 199.28 0.46 ;
    RECT 197.01 0.0 197.72 0.46 ;
    RECT 195.99 0.0 196.49 0.46 ;
    RECT 193.6 0.0 194.1 0.46 ;
    RECT 192.37 0.0 193.08 0.46 ;
    RECT 190.81 0.0 191.52 0.46 ;
    RECT 189.79 0.0 190.29 0.46 ;
    RECT 187.4 0.0 187.9 0.46 ;
    RECT 186.17 0.0 186.88 0.46 ;
    RECT 184.61 0.0 185.32 0.46 ;
    RECT 183.59 0.0 184.09 0.46 ;
    RECT 181.2 0.0 181.7 0.46 ;
    RECT 179.97 0.0 180.68 0.46 ;
    RECT 178.41 0.0 179.12 0.46 ;
    RECT 177.39 0.0 177.89 0.46 ;
    RECT 175.0 0.0 175.5 0.46 ;
    RECT 173.77 0.0 174.48 0.46 ;
    RECT 172.21 0.0 172.92 0.46 ;
    RECT 171.19 0.0 171.69 0.46 ;
    RECT 168.8 0.0 169.3 0.46 ;
    RECT 167.57 0.0 168.28 0.46 ;
    RECT 166.01 0.0 166.72 0.46 ;
    RECT 164.99 0.0 165.49 0.46 ;
    RECT 162.815 0.0 163.94 0.46 ;
    RECT 162.425 0.0 162.605 0.46 ;
    RECT 160.545 0.0 162.215 0.46 ;
    RECT 159.48 0.0 160.335 0.46 ;
    RECT 156.82 0.0 159.27 0.46 ;
    RECT 156.5 0.0 156.61 0.46 ;
    RECT 154.835 0.0 156.29 0.46 ;
    RECT 154.515 0.0 154.625 0.46 ;
    RECT 152.71 0.0 154.305 0.46 ;
    RECT 151.375 0.0 152.5 0.46 ;
    RECT 151.055 0.0 151.165 0.46 ;
    RECT 150.355 0.0 150.845 0.46 ;
    RECT 149.465 0.0 150.145 0.46 ;
    RECT 148.405 0.0 149.255 0.46 ;
    RECT 148.085 0.0 148.195 0.46 ;
    RECT 147.175 0.0 147.875 0.46 ;
    RECT 145.14 0.0 146.965 0.46 ;
    RECT 143.95 0.0 144.93 0.46 ;
    RECT 141.915 0.0 143.74 0.46 ;
    RECT 141.005 0.0 141.705 0.46 ;
    RECT 140.685 0.0 140.795 0.46 ;
    RECT 139.625 0.0 140.475 0.46 ;
    RECT 138.735 0.0 139.415 0.46 ;
    RECT 138.035 0.0 138.525 0.46 ;
    RECT 137.715 0.0 137.825 0.46 ;
    RECT 136.66 0.0 137.505 0.46 ;
    RECT 134.575 0.0 136.17 0.46 ;
    RECT 134.255 0.0 134.365 0.46 ;
    RECT 132.59 0.0 134.045 0.46 ;
    RECT 132.27 0.0 132.38 0.46 ;
    RECT 129.61 0.0 132.06 0.46 ;
    RECT 128.545 0.0 129.4 0.46 ;
    RECT 126.665 0.0 128.335 0.46 ;
    RECT 126.275 0.0 126.455 0.46 ;
    RECT 124.94 0.0 126.065 0.46 ;
    RECT 123.39 0.0 123.89 0.46 ;
    RECT 122.16 0.0 122.87 0.46 ;
    RECT 120.6 0.0 121.31 0.46 ;
    RECT 119.58 0.0 120.08 0.46 ;
    RECT 117.19 0.0 117.69 0.46 ;
    RECT 115.96 0.0 116.67 0.46 ;
    RECT 114.4 0.0 115.11 0.46 ;
    RECT 113.38 0.0 113.88 0.46 ;
    RECT 110.99 0.0 111.49 0.46 ;
    RECT 109.76 0.0 110.47 0.46 ;
    RECT 108.2 0.0 108.91 0.46 ;
    RECT 107.18 0.0 107.68 0.46 ;
    RECT 104.79 0.0 105.29 0.46 ;
    RECT 103.56 0.0 104.27 0.46 ;
    RECT 102.0 0.0 102.71 0.46 ;
    RECT 100.98 0.0 101.48 0.46 ;
    RECT 98.59 0.0 99.09 0.46 ;
    RECT 97.36 0.0 98.07 0.46 ;
    RECT 95.8 0.0 96.51 0.46 ;
    RECT 94.78 0.0 95.28 0.46 ;
    RECT 92.39 0.0 92.89 0.46 ;
    RECT 91.16 0.0 91.87 0.46 ;
    RECT 89.6 0.0 90.31 0.46 ;
    RECT 88.58 0.0 89.08 0.46 ;
    RECT 86.19 0.0 86.69 0.46 ;
    RECT 84.96 0.0 85.67 0.46 ;
    RECT 83.4 0.0 84.11 0.46 ;
    RECT 82.38 0.0 82.88 0.46 ;
    RECT 79.99 0.0 80.49 0.46 ;
    RECT 78.76 0.0 79.47 0.46 ;
    RECT 77.2 0.0 77.91 0.46 ;
    RECT 76.18 0.0 76.68 0.46 ;
    RECT 73.79 0.0 74.29 0.46 ;
    RECT 72.56 0.0 73.27 0.46 ;
    RECT 71.0 0.0 71.71 0.46 ;
    RECT 69.98 0.0 70.48 0.46 ;
    RECT 67.59 0.0 68.09 0.46 ;
    RECT 66.36 0.0 67.07 0.46 ;
    RECT 64.8 0.0 65.51 0.46 ;
    RECT 63.78 0.0 64.28 0.46 ;
    RECT 61.39 0.0 61.89 0.46 ;
    RECT 60.16 0.0 60.87 0.46 ;
    RECT 58.6 0.0 59.31 0.46 ;
    RECT 57.58 0.0 58.08 0.46 ;
    RECT 55.19 0.0 55.69 0.46 ;
    RECT 53.96 0.0 54.67 0.46 ;
    RECT 52.4 0.0 53.11 0.46 ;
    RECT 51.38 0.0 51.88 0.46 ;
    RECT 48.99 0.0 49.49 0.46 ;
    RECT 47.76 0.0 48.47 0.46 ;
    RECT 46.2 0.0 46.91 0.46 ;
    RECT 45.18 0.0 45.68 0.46 ;
    RECT 42.79 0.0 43.29 0.46 ;
    RECT 41.56 0.0 42.27 0.46 ;
    RECT 40.0 0.0 40.71 0.46 ;
    RECT 38.98 0.0 39.48 0.46 ;
    RECT 36.59 0.0 37.09 0.46 ;
    RECT 35.36 0.0 36.07 0.46 ;
    RECT 33.8 0.0 34.51 0.46 ;
    RECT 32.78 0.0 33.28 0.46 ;
    RECT 30.39 0.0 30.89 0.46 ;
    RECT 29.16 0.0 29.87 0.46 ;
    RECT 27.6 0.0 28.31 0.46 ;
    RECT 26.58 0.0 27.08 0.46 ;
    RECT 24.19 0.0 24.69 0.46 ;
    RECT 22.96 0.0 23.67 0.46 ;
    RECT 21.4 0.0 22.11 0.46 ;
    RECT 20.38 0.0 20.88 0.46 ;
    RECT 17.99 0.0 18.49 0.46 ;
    RECT 16.76 0.0 17.47 0.46 ;
    RECT 15.2 0.0 15.91 0.46 ;
    RECT 14.18 0.0 14.68 0.46 ;
    RECT 11.79 0.0 12.29 0.46 ;
    RECT 10.56 0.0 11.27 0.46 ;
    RECT 9.0 0.0 9.71 0.46 ;
    RECT 7.98 0.0 8.48 0.46 ;
    RECT 5.59 0.0 6.09 0.46 ;
    RECT 4.36 0.0 5.07 0.46 ;
    RECT 2.8 0.0 3.51 0.46 ;
    RECT 1.78 0.0 2.28 0.46 ;
    RECT 0.59 0.0 0.73 0.46 ;
    RECT 0.0 0.0 0.38 0.46 ;
    RECT 576.8 0.46 577.18 270.08 ;
    RECT 576.45 0.46 576.59 270.08 ;
    RECT 575.61 0.46 576.24 270.08 ;
    RECT 574.9 0.46 575.4 270.08 ;
    RECT 573.35 0.46 574.69 270.08 ;
    RECT 571.8 0.46 573.14 270.08 ;
    RECT 571.09 0.46 571.59 270.08 ;
    RECT 570.25 0.46 570.88 270.08 ;
    RECT 569.41 0.46 570.04 270.08 ;
    RECT 568.7 0.46 569.2 270.08 ;
    RECT 567.15 0.46 568.49 270.08 ;
    RECT 565.6 0.46 566.94 270.08 ;
    RECT 564.89 0.46 565.39 270.08 ;
    RECT 564.05 0.46 564.68 270.08 ;
    RECT 563.21 0.46 563.84 270.08 ;
    RECT 562.5 0.46 563.0 270.08 ;
    RECT 560.95 0.46 562.29 270.08 ;
    RECT 559.4 0.46 560.74 270.08 ;
    RECT 558.69 0.46 559.19 270.08 ;
    RECT 557.85 0.46 558.48 270.08 ;
    RECT 557.01 0.46 557.64 270.08 ;
    RECT 556.3 0.46 556.8 270.08 ;
    RECT 554.75 0.46 556.09 270.08 ;
    RECT 553.2 0.46 554.54 270.08 ;
    RECT 552.49 0.46 552.99 270.08 ;
    RECT 551.65 0.46 552.28 270.08 ;
    RECT 550.81 0.46 551.44 270.08 ;
    RECT 550.1 0.46 550.6 270.08 ;
    RECT 548.55 0.46 549.89 270.08 ;
    RECT 547.0 0.46 548.34 270.08 ;
    RECT 546.29 0.46 546.79 270.08 ;
    RECT 545.45 0.46 546.08 270.08 ;
    RECT 544.61 0.46 545.24 270.08 ;
    RECT 543.9 0.46 544.4 270.08 ;
    RECT 542.35 0.46 543.69 270.08 ;
    RECT 540.8 0.46 542.14 270.08 ;
    RECT 540.09 0.46 540.59 270.08 ;
    RECT 539.25 0.46 539.88 270.08 ;
    RECT 538.41 0.46 539.04 270.08 ;
    RECT 537.7 0.46 538.2 270.08 ;
    RECT 536.15 0.46 537.49 270.08 ;
    RECT 534.6 0.46 535.94 270.08 ;
    RECT 533.89 0.46 534.39 270.08 ;
    RECT 533.05 0.46 533.68 270.08 ;
    RECT 532.21 0.46 532.84 270.08 ;
    RECT 531.5 0.46 532.0 270.08 ;
    RECT 529.95 0.46 531.29 270.08 ;
    RECT 528.4 0.46 529.74 270.08 ;
    RECT 527.69 0.46 528.19 270.08 ;
    RECT 526.85 0.46 527.48 270.08 ;
    RECT 526.01 0.46 526.64 270.08 ;
    RECT 525.3 0.46 525.8 270.08 ;
    RECT 523.75 0.46 525.09 270.08 ;
    RECT 522.2 0.46 523.54 270.08 ;
    RECT 521.49 0.46 521.99 270.08 ;
    RECT 520.65 0.46 521.28 270.08 ;
    RECT 519.81 0.46 520.44 270.08 ;
    RECT 519.1 0.46 519.6 270.08 ;
    RECT 517.55 0.46 518.89 270.08 ;
    RECT 516.0 0.46 517.34 270.08 ;
    RECT 515.29 0.46 515.79 270.08 ;
    RECT 514.45 0.46 515.08 270.08 ;
    RECT 513.61 0.46 514.24 270.08 ;
    RECT 512.9 0.46 513.4 270.08 ;
    RECT 511.35 0.46 512.69 270.08 ;
    RECT 509.8 0.46 511.14 270.08 ;
    RECT 509.09 0.46 509.59 270.08 ;
    RECT 508.25 0.46 508.88 270.08 ;
    RECT 507.41 0.46 508.04 270.08 ;
    RECT 506.7 0.46 507.2 270.08 ;
    RECT 505.15 0.46 506.49 270.08 ;
    RECT 503.6 0.46 504.94 270.08 ;
    RECT 502.89 0.46 503.39 270.08 ;
    RECT 502.05 0.46 502.68 270.08 ;
    RECT 501.21 0.46 501.84 270.08 ;
    RECT 500.5 0.46 501.0 270.08 ;
    RECT 498.95 0.46 500.29 270.08 ;
    RECT 497.4 0.46 498.74 270.08 ;
    RECT 496.69 0.46 497.19 270.08 ;
    RECT 495.85 0.46 496.48 270.08 ;
    RECT 495.01 0.46 495.64 270.08 ;
    RECT 494.3 0.46 494.8 270.08 ;
    RECT 492.75 0.46 494.09 270.08 ;
    RECT 491.2 0.46 492.54 270.08 ;
    RECT 490.49 0.46 490.99 270.08 ;
    RECT 489.65 0.46 490.28 270.08 ;
    RECT 488.81 0.46 489.44 270.08 ;
    RECT 488.1 0.46 488.6 270.08 ;
    RECT 486.55 0.46 487.89 270.08 ;
    RECT 485.0 0.46 486.34 270.08 ;
    RECT 484.29 0.46 484.79 270.08 ;
    RECT 483.45 0.46 484.08 270.08 ;
    RECT 482.61 0.46 483.24 270.08 ;
    RECT 481.9 0.46 482.4 270.08 ;
    RECT 480.35 0.46 481.69 270.08 ;
    RECT 478.8 0.46 480.14 270.08 ;
    RECT 478.09 0.46 478.59 270.08 ;
    RECT 477.25 0.46 477.88 270.08 ;
    RECT 476.41 0.46 477.04 270.08 ;
    RECT 475.7 0.46 476.2 270.08 ;
    RECT 474.15 0.46 475.49 270.08 ;
    RECT 472.6 0.46 473.94 270.08 ;
    RECT 471.89 0.46 472.39 270.08 ;
    RECT 471.05 0.46 471.68 270.08 ;
    RECT 470.21 0.46 470.84 270.08 ;
    RECT 469.5 0.46 470.0 270.08 ;
    RECT 467.95 0.46 469.29 270.08 ;
    RECT 466.4 0.46 467.74 270.08 ;
    RECT 465.69 0.46 466.19 270.08 ;
    RECT 464.85 0.46 465.48 270.08 ;
    RECT 464.01 0.46 464.64 270.08 ;
    RECT 463.3 0.46 463.8 270.08 ;
    RECT 461.75 0.46 463.09 270.08 ;
    RECT 460.2 0.46 461.54 270.08 ;
    RECT 459.49 0.46 459.99 270.08 ;
    RECT 458.65 0.46 459.28 270.08 ;
    RECT 457.81 0.46 458.44 270.08 ;
    RECT 457.1 0.46 457.6 270.08 ;
    RECT 455.55 0.46 456.89 270.08 ;
    RECT 454.0 0.46 455.34 270.08 ;
    RECT 453.29 0.46 453.79 270.08 ;
    RECT 452.45 0.46 453.08 270.08 ;
    RECT 451.115 0.46 452.24 270.08 ;
    RECT 450.725 0.46 450.905 270.08 ;
    RECT 448.845 0.46 450.515 270.08 ;
    RECT 447.78 0.46 448.635 270.08 ;
    RECT 445.12 0.46 447.57 270.08 ;
    RECT 444.8 0.46 444.91 270.08 ;
    RECT 443.135 0.46 444.59 270.08 ;
    RECT 442.815 0.46 442.925 270.08 ;
    RECT 441.01 0.46 442.605 270.08 ;
    RECT 439.675 0.46 440.52 270.08 ;
    RECT 439.355 0.46 439.465 270.08 ;
    RECT 438.655 0.46 439.145 270.08 ;
    RECT 437.765 0.46 438.445 270.08 ;
    RECT 436.705 0.46 437.555 270.08 ;
    RECT 436.385 0.46 436.495 270.08 ;
    RECT 435.475 0.46 436.175 270.08 ;
    RECT 433.44 0.46 435.265 270.08 ;
    RECT 432.25 0.46 433.23 270.08 ;
    RECT 430.215 0.46 432.04 270.08 ;
    RECT 429.305 0.46 430.005 270.08 ;
    RECT 428.985 0.46 429.095 270.08 ;
    RECT 427.925 0.46 428.775 270.08 ;
    RECT 427.035 0.46 427.715 270.08 ;
    RECT 426.335 0.46 426.825 270.08 ;
    RECT 426.015 0.46 426.125 270.08 ;
    RECT 424.68 0.46 425.805 270.08 ;
    RECT 422.875 0.46 424.47 270.08 ;
    RECT 422.555 0.46 422.665 270.08 ;
    RECT 420.89 0.46 422.345 270.08 ;
    RECT 420.57 0.46 420.68 270.08 ;
    RECT 417.91 0.46 420.36 270.08 ;
    RECT 416.845 0.46 417.7 270.08 ;
    RECT 414.965 0.46 416.635 270.08 ;
    RECT 414.575 0.46 414.755 270.08 ;
    RECT 413.24 0.46 414.365 270.08 ;
    RECT 412.4 0.46 413.03 270.08 ;
    RECT 411.69 0.46 412.19 270.08 ;
    RECT 410.14 0.46 411.48 270.08 ;
    RECT 408.59 0.46 409.93 270.08 ;
    RECT 407.88 0.46 408.38 270.08 ;
    RECT 407.04 0.46 407.67 270.08 ;
    RECT 406.2 0.46 406.83 270.08 ;
    RECT 405.49 0.46 405.99 270.08 ;
    RECT 403.94 0.46 405.28 270.08 ;
    RECT 402.39 0.46 403.73 270.08 ;
    RECT 401.68 0.46 402.18 270.08 ;
    RECT 400.84 0.46 401.47 270.08 ;
    RECT 400.0 0.46 400.63 270.08 ;
    RECT 399.29 0.46 399.79 270.08 ;
    RECT 397.74 0.46 399.08 270.08 ;
    RECT 396.19 0.46 397.53 270.08 ;
    RECT 395.48 0.46 395.98 270.08 ;
    RECT 394.64 0.46 395.27 270.08 ;
    RECT 393.8 0.46 394.43 270.08 ;
    RECT 393.09 0.46 393.59 270.08 ;
    RECT 391.54 0.46 392.88 270.08 ;
    RECT 389.99 0.46 391.33 270.08 ;
    RECT 389.28 0.46 389.78 270.08 ;
    RECT 388.44 0.46 389.07 270.08 ;
    RECT 387.6 0.46 388.23 270.08 ;
    RECT 386.89 0.46 387.39 270.08 ;
    RECT 385.34 0.46 386.68 270.08 ;
    RECT 383.79 0.46 385.13 270.08 ;
    RECT 383.08 0.46 383.58 270.08 ;
    RECT 382.24 0.46 382.87 270.08 ;
    RECT 381.4 0.46 382.03 270.08 ;
    RECT 380.69 0.46 381.19 270.08 ;
    RECT 379.14 0.46 380.48 270.08 ;
    RECT 377.59 0.46 378.93 270.08 ;
    RECT 376.88 0.46 377.38 270.08 ;
    RECT 376.04 0.46 376.67 270.08 ;
    RECT 375.2 0.46 375.83 270.08 ;
    RECT 374.49 0.46 374.99 270.08 ;
    RECT 372.94 0.46 374.28 270.08 ;
    RECT 371.39 0.46 372.73 270.08 ;
    RECT 370.68 0.46 371.18 270.08 ;
    RECT 369.84 0.46 370.47 270.08 ;
    RECT 369.0 0.46 369.63 270.08 ;
    RECT 368.29 0.46 368.79 270.08 ;
    RECT 366.74 0.46 368.08 270.08 ;
    RECT 365.19 0.46 366.53 270.08 ;
    RECT 364.48 0.46 364.98 270.08 ;
    RECT 363.64 0.46 364.27 270.08 ;
    RECT 362.8 0.46 363.43 270.08 ;
    RECT 362.09 0.46 362.59 270.08 ;
    RECT 360.54 0.46 361.88 270.08 ;
    RECT 358.99 0.46 360.33 270.08 ;
    RECT 358.28 0.46 358.78 270.08 ;
    RECT 357.44 0.46 358.07 270.08 ;
    RECT 356.6 0.46 357.23 270.08 ;
    RECT 355.89 0.46 356.39 270.08 ;
    RECT 354.34 0.46 355.68 270.08 ;
    RECT 352.79 0.46 354.13 270.08 ;
    RECT 352.08 0.46 352.58 270.08 ;
    RECT 351.24 0.46 351.87 270.08 ;
    RECT 350.4 0.46 351.03 270.08 ;
    RECT 349.69 0.46 350.19 270.08 ;
    RECT 348.14 0.46 349.48 270.08 ;
    RECT 346.59 0.46 347.93 270.08 ;
    RECT 345.88 0.46 346.38 270.08 ;
    RECT 345.04 0.46 345.67 270.08 ;
    RECT 344.2 0.46 344.83 270.08 ;
    RECT 343.49 0.46 343.99 270.08 ;
    RECT 341.94 0.46 343.28 270.08 ;
    RECT 340.39 0.46 341.73 270.08 ;
    RECT 339.68 0.46 340.18 270.08 ;
    RECT 338.84 0.46 339.47 270.08 ;
    RECT 338.0 0.46 338.63 270.08 ;
    RECT 337.29 0.46 337.79 270.08 ;
    RECT 335.74 0.46 337.08 270.08 ;
    RECT 334.19 0.46 335.53 270.08 ;
    RECT 333.48 0.46 333.98 270.08 ;
    RECT 332.64 0.46 333.27 270.08 ;
    RECT 331.8 0.46 332.43 270.08 ;
    RECT 331.09 0.46 331.59 270.08 ;
    RECT 329.54 0.46 330.88 270.08 ;
    RECT 327.99 0.46 329.33 270.08 ;
    RECT 327.28 0.46 327.78 270.08 ;
    RECT 326.44 0.46 327.07 270.08 ;
    RECT 325.6 0.46 326.23 270.08 ;
    RECT 324.89 0.46 325.39 270.08 ;
    RECT 323.34 0.46 324.68 270.08 ;
    RECT 321.79 0.46 323.13 270.08 ;
    RECT 321.08 0.46 321.58 270.08 ;
    RECT 320.24 0.46 320.87 270.08 ;
    RECT 319.4 0.46 320.03 270.08 ;
    RECT 318.69 0.46 319.19 270.08 ;
    RECT 317.14 0.46 318.48 270.08 ;
    RECT 315.59 0.46 316.93 270.08 ;
    RECT 314.88 0.46 315.38 270.08 ;
    RECT 314.04 0.46 314.67 270.08 ;
    RECT 313.2 0.46 313.83 270.08 ;
    RECT 312.49 0.46 312.99 270.08 ;
    RECT 310.94 0.46 312.28 270.08 ;
    RECT 309.39 0.46 310.73 270.08 ;
    RECT 308.68 0.46 309.18 270.08 ;
    RECT 307.84 0.46 308.47 270.08 ;
    RECT 307.0 0.46 307.63 270.08 ;
    RECT 306.29 0.46 306.79 270.08 ;
    RECT 304.74 0.46 306.08 270.08 ;
    RECT 303.19 0.46 304.53 270.08 ;
    RECT 302.48 0.46 302.98 270.08 ;
    RECT 301.64 0.46 302.27 270.08 ;
    RECT 300.8 0.46 301.43 270.08 ;
    RECT 300.09 0.46 300.59 270.08 ;
    RECT 298.54 0.46 299.88 270.08 ;
    RECT 296.99 0.46 298.33 270.08 ;
    RECT 296.28 0.46 296.78 270.08 ;
    RECT 295.44 0.46 296.07 270.08 ;
    RECT 294.6 0.46 295.23 270.08 ;
    RECT 293.89 0.46 294.39 270.08 ;
    RECT 292.34 0.46 293.68 270.08 ;
    RECT 290.79 0.46 292.13 270.08 ;
    RECT 290.08 0.46 290.58 270.08 ;
    RECT 289.24 0.46 289.87 270.08 ;
    RECT 288.15 0.46 289.03 270.08 ;
    RECT 287.31 0.46 287.94 270.08 ;
    RECT 286.6 0.46 287.1 270.08 ;
    RECT 285.05 0.46 286.39 270.08 ;
    RECT 283.5 0.46 284.84 270.08 ;
    RECT 282.79 0.46 283.29 270.08 ;
    RECT 281.95 0.46 282.58 270.08 ;
    RECT 281.11 0.46 281.74 270.08 ;
    RECT 280.4 0.46 280.9 270.08 ;
    RECT 278.85 0.46 280.19 270.08 ;
    RECT 277.3 0.46 278.64 270.08 ;
    RECT 276.59 0.46 277.09 270.08 ;
    RECT 275.75 0.46 276.38 270.08 ;
    RECT 274.91 0.46 275.54 270.08 ;
    RECT 274.2 0.46 274.7 270.08 ;
    RECT 272.65 0.46 273.99 270.08 ;
    RECT 271.1 0.46 272.44 270.08 ;
    RECT 270.39 0.46 270.89 270.08 ;
    RECT 269.55 0.46 270.18 270.08 ;
    RECT 268.71 0.46 269.34 270.08 ;
    RECT 268.0 0.46 268.5 270.08 ;
    RECT 266.45 0.46 267.79 270.08 ;
    RECT 264.9 0.46 266.24 270.08 ;
    RECT 264.19 0.46 264.69 270.08 ;
    RECT 263.35 0.46 263.98 270.08 ;
    RECT 262.51 0.46 263.14 270.08 ;
    RECT 261.8 0.46 262.3 270.08 ;
    RECT 260.25 0.46 261.59 270.08 ;
    RECT 258.7 0.46 260.04 270.08 ;
    RECT 257.99 0.46 258.49 270.08 ;
    RECT 257.15 0.46 257.78 270.08 ;
    RECT 256.31 0.46 256.94 270.08 ;
    RECT 255.6 0.46 256.1 270.08 ;
    RECT 254.05 0.46 255.39 270.08 ;
    RECT 252.5 0.46 253.84 270.08 ;
    RECT 251.79 0.46 252.29 270.08 ;
    RECT 250.95 0.46 251.58 270.08 ;
    RECT 250.11 0.46 250.74 270.08 ;
    RECT 249.4 0.46 249.9 270.08 ;
    RECT 247.85 0.46 249.19 270.08 ;
    RECT 246.3 0.46 247.64 270.08 ;
    RECT 245.59 0.46 246.09 270.08 ;
    RECT 244.75 0.46 245.38 270.08 ;
    RECT 243.91 0.46 244.54 270.08 ;
    RECT 243.2 0.46 243.7 270.08 ;
    RECT 241.65 0.46 242.99 270.08 ;
    RECT 240.1 0.46 241.44 270.08 ;
    RECT 239.39 0.46 239.89 270.08 ;
    RECT 238.55 0.46 239.18 270.08 ;
    RECT 237.71 0.46 238.34 270.08 ;
    RECT 237.0 0.46 237.5 270.08 ;
    RECT 235.45 0.46 236.79 270.08 ;
    RECT 233.9 0.46 235.24 270.08 ;
    RECT 233.19 0.46 233.69 270.08 ;
    RECT 232.35 0.46 232.98 270.08 ;
    RECT 231.51 0.46 232.14 270.08 ;
    RECT 230.8 0.46 231.3 270.08 ;
    RECT 229.25 0.46 230.59 270.08 ;
    RECT 227.7 0.46 229.04 270.08 ;
    RECT 226.99 0.46 227.49 270.08 ;
    RECT 226.15 0.46 226.78 270.08 ;
    RECT 225.31 0.46 225.94 270.08 ;
    RECT 224.6 0.46 225.1 270.08 ;
    RECT 223.05 0.46 224.39 270.08 ;
    RECT 221.5 0.46 222.84 270.08 ;
    RECT 220.79 0.46 221.29 270.08 ;
    RECT 219.95 0.46 220.58 270.08 ;
    RECT 219.11 0.46 219.74 270.08 ;
    RECT 218.4 0.46 218.9 270.08 ;
    RECT 216.85 0.46 218.19 270.08 ;
    RECT 215.3 0.46 216.64 270.08 ;
    RECT 214.59 0.46 215.09 270.08 ;
    RECT 213.75 0.46 214.38 270.08 ;
    RECT 212.91 0.46 213.54 270.08 ;
    RECT 212.2 0.46 212.7 270.08 ;
    RECT 210.65 0.46 211.99 270.08 ;
    RECT 209.1 0.46 210.44 270.08 ;
    RECT 208.39 0.46 208.89 270.08 ;
    RECT 207.55 0.46 208.18 270.08 ;
    RECT 206.71 0.46 207.34 270.08 ;
    RECT 206.0 0.46 206.5 270.08 ;
    RECT 204.45 0.46 205.79 270.08 ;
    RECT 202.9 0.46 204.24 270.08 ;
    RECT 202.19 0.46 202.69 270.08 ;
    RECT 201.35 0.46 201.98 270.08 ;
    RECT 200.51 0.46 201.14 270.08 ;
    RECT 199.8 0.46 200.3 270.08 ;
    RECT 198.25 0.46 199.59 270.08 ;
    RECT 196.7 0.46 198.04 270.08 ;
    RECT 195.99 0.46 196.49 270.08 ;
    RECT 195.15 0.46 195.78 270.08 ;
    RECT 194.31 0.46 194.94 270.08 ;
    RECT 193.6 0.46 194.1 270.08 ;
    RECT 192.05 0.46 193.39 270.08 ;
    RECT 190.5 0.46 191.84 270.08 ;
    RECT 189.79 0.46 190.29 270.08 ;
    RECT 188.95 0.46 189.58 270.08 ;
    RECT 188.11 0.46 188.74 270.08 ;
    RECT 187.4 0.46 187.9 270.08 ;
    RECT 185.85 0.46 187.19 270.08 ;
    RECT 184.3 0.46 185.64 270.08 ;
    RECT 183.59 0.46 184.09 270.08 ;
    RECT 182.75 0.46 183.38 270.08 ;
    RECT 181.91 0.46 182.54 270.08 ;
    RECT 181.2 0.46 181.7 270.08 ;
    RECT 179.65 0.46 180.99 270.08 ;
    RECT 178.1 0.46 179.44 270.08 ;
    RECT 177.39 0.46 177.89 270.08 ;
    RECT 176.55 0.46 177.18 270.08 ;
    RECT 175.71 0.46 176.34 270.08 ;
    RECT 175.0 0.46 175.5 270.08 ;
    RECT 173.45 0.46 174.79 270.08 ;
    RECT 171.9 0.46 173.24 270.08 ;
    RECT 171.19 0.46 171.69 270.08 ;
    RECT 170.35 0.46 170.98 270.08 ;
    RECT 169.51 0.46 170.14 270.08 ;
    RECT 168.8 0.46 169.3 270.08 ;
    RECT 167.25 0.46 168.59 270.08 ;
    RECT 165.7 0.46 167.04 270.08 ;
    RECT 164.99 0.46 165.49 270.08 ;
    RECT 164.15 0.46 164.78 270.08 ;
    RECT 162.815 0.46 163.94 270.08 ;
    RECT 162.425 0.46 162.605 270.08 ;
    RECT 160.545 0.46 162.215 270.08 ;
    RECT 159.48 0.46 160.335 270.08 ;
    RECT 156.82 0.46 159.27 270.08 ;
    RECT 156.5 0.46 156.61 270.08 ;
    RECT 154.835 0.46 156.29 270.08 ;
    RECT 154.515 0.46 154.625 270.08 ;
    RECT 152.71 0.46 154.305 270.08 ;
    RECT 151.375 0.46 152.5 270.08 ;
    RECT 151.055 0.46 151.165 270.08 ;
    RECT 150.355 0.46 150.845 270.08 ;
    RECT 149.465 0.46 150.145 270.08 ;
    RECT 148.405 0.46 149.255 270.08 ;
    RECT 148.085 0.46 148.195 270.08 ;
    RECT 147.175 0.46 147.875 270.08 ;
    RECT 145.14 0.46 146.965 270.08 ;
    RECT 143.95 0.46 144.93 270.08 ;
    RECT 141.915 0.46 143.74 270.08 ;
    RECT 141.005 0.46 141.705 270.08 ;
    RECT 140.685 0.46 140.795 270.08 ;
    RECT 139.625 0.46 140.475 270.08 ;
    RECT 138.735 0.46 139.415 270.08 ;
    RECT 138.035 0.46 138.525 270.08 ;
    RECT 137.715 0.46 137.825 270.08 ;
    RECT 136.66 0.46 137.505 270.08 ;
    RECT 134.575 0.46 136.17 270.08 ;
    RECT 134.255 0.46 134.365 270.08 ;
    RECT 132.59 0.46 134.045 270.08 ;
    RECT 132.27 0.46 132.38 270.08 ;
    RECT 129.61 0.46 132.06 270.08 ;
    RECT 128.545 0.46 129.4 270.08 ;
    RECT 126.665 0.46 128.335 270.08 ;
    RECT 126.275 0.46 126.455 270.08 ;
    RECT 124.94 0.46 126.065 270.08 ;
    RECT 124.1 0.46 124.73 270.08 ;
    RECT 123.39 0.46 123.89 270.08 ;
    RECT 121.84 0.46 123.18 270.08 ;
    RECT 120.29 0.46 121.63 270.08 ;
    RECT 119.58 0.46 120.08 270.08 ;
    RECT 118.74 0.46 119.37 270.08 ;
    RECT 117.9 0.46 118.53 270.08 ;
    RECT 117.19 0.46 117.69 270.08 ;
    RECT 115.64 0.46 116.98 270.08 ;
    RECT 114.09 0.46 115.43 270.08 ;
    RECT 113.38 0.46 113.88 270.08 ;
    RECT 112.54 0.46 113.17 270.08 ;
    RECT 111.7 0.46 112.33 270.08 ;
    RECT 110.99 0.46 111.49 270.08 ;
    RECT 109.44 0.46 110.78 270.08 ;
    RECT 107.89 0.46 109.23 270.08 ;
    RECT 107.18 0.46 107.68 270.08 ;
    RECT 106.34 0.46 106.97 270.08 ;
    RECT 105.5 0.46 106.13 270.08 ;
    RECT 104.79 0.46 105.29 270.08 ;
    RECT 103.24 0.46 104.58 270.08 ;
    RECT 101.69 0.46 103.03 270.08 ;
    RECT 100.98 0.46 101.48 270.08 ;
    RECT 100.14 0.46 100.77 270.08 ;
    RECT 99.3 0.46 99.93 270.08 ;
    RECT 98.59 0.46 99.09 270.08 ;
    RECT 97.04 0.46 98.38 270.08 ;
    RECT 95.49 0.46 96.83 270.08 ;
    RECT 94.78 0.46 95.28 270.08 ;
    RECT 93.94 0.46 94.57 270.08 ;
    RECT 93.1 0.46 93.73 270.08 ;
    RECT 92.39 0.46 92.89 270.08 ;
    RECT 90.84 0.46 92.18 270.08 ;
    RECT 89.29 0.46 90.63 270.08 ;
    RECT 88.58 0.46 89.08 270.08 ;
    RECT 87.74 0.46 88.37 270.08 ;
    RECT 86.9 0.46 87.53 270.08 ;
    RECT 86.19 0.46 86.69 270.08 ;
    RECT 84.64 0.46 85.98 270.08 ;
    RECT 83.09 0.46 84.43 270.08 ;
    RECT 82.38 0.46 82.88 270.08 ;
    RECT 81.54 0.46 82.17 270.08 ;
    RECT 80.7 0.46 81.33 270.08 ;
    RECT 79.99 0.46 80.49 270.08 ;
    RECT 78.44 0.46 79.78 270.08 ;
    RECT 76.89 0.46 78.23 270.08 ;
    RECT 76.18 0.46 76.68 270.08 ;
    RECT 75.34 0.46 75.97 270.08 ;
    RECT 74.5 0.46 75.13 270.08 ;
    RECT 73.79 0.46 74.29 270.08 ;
    RECT 72.24 0.46 73.58 270.08 ;
    RECT 70.69 0.46 72.03 270.08 ;
    RECT 69.98 0.46 70.48 270.08 ;
    RECT 69.14 0.46 69.77 270.08 ;
    RECT 68.3 0.46 68.93 270.08 ;
    RECT 67.59 0.46 68.09 270.08 ;
    RECT 66.04 0.46 67.38 270.08 ;
    RECT 64.49 0.46 65.83 270.08 ;
    RECT 63.78 0.46 64.28 270.08 ;
    RECT 62.94 0.46 63.57 270.08 ;
    RECT 62.1 0.46 62.73 270.08 ;
    RECT 61.39 0.46 61.89 270.08 ;
    RECT 59.84 0.46 61.18 270.08 ;
    RECT 58.29 0.46 59.63 270.08 ;
    RECT 57.58 0.46 58.08 270.08 ;
    RECT 56.74 0.46 57.37 270.08 ;
    RECT 55.9 0.46 56.53 270.08 ;
    RECT 55.19 0.46 55.69 270.08 ;
    RECT 53.64 0.46 54.98 270.08 ;
    RECT 52.09 0.46 53.43 270.08 ;
    RECT 51.38 0.46 51.88 270.08 ;
    RECT 50.54 0.46 51.17 270.08 ;
    RECT 49.7 0.46 50.33 270.08 ;
    RECT 48.99 0.46 49.49 270.08 ;
    RECT 47.44 0.46 48.78 270.08 ;
    RECT 45.89 0.46 47.23 270.08 ;
    RECT 45.18 0.46 45.68 270.08 ;
    RECT 44.34 0.46 44.97 270.08 ;
    RECT 43.5 0.46 44.13 270.08 ;
    RECT 42.79 0.46 43.29 270.08 ;
    RECT 41.24 0.46 42.58 270.08 ;
    RECT 39.69 0.46 41.03 270.08 ;
    RECT 38.98 0.46 39.48 270.08 ;
    RECT 38.14 0.46 38.77 270.08 ;
    RECT 37.3 0.46 37.93 270.08 ;
    RECT 36.59 0.46 37.09 270.08 ;
    RECT 35.04 0.46 36.38 270.08 ;
    RECT 33.49 0.46 34.83 270.08 ;
    RECT 32.78 0.46 33.28 270.08 ;
    RECT 31.94 0.46 32.57 270.08 ;
    RECT 31.1 0.46 31.73 270.08 ;
    RECT 30.39 0.46 30.89 270.08 ;
    RECT 28.84 0.46 30.18 270.08 ;
    RECT 27.29 0.46 28.63 270.08 ;
    RECT 26.58 0.46 27.08 270.08 ;
    RECT 25.74 0.46 26.37 270.08 ;
    RECT 24.9 0.46 25.53 270.08 ;
    RECT 24.19 0.46 24.69 270.08 ;
    RECT 22.64 0.46 23.98 270.08 ;
    RECT 21.09 0.46 22.43 270.08 ;
    RECT 20.38 0.46 20.88 270.08 ;
    RECT 19.54 0.46 20.17 270.08 ;
    RECT 18.7 0.46 19.33 270.08 ;
    RECT 17.99 0.46 18.49 270.08 ;
    RECT 16.44 0.46 17.78 270.08 ;
    RECT 14.89 0.46 16.23 270.08 ;
    RECT 14.18 0.46 14.68 270.08 ;
    RECT 13.34 0.46 13.97 270.08 ;
    RECT 12.5 0.46 13.13 270.08 ;
    RECT 11.79 0.46 12.29 270.08 ;
    RECT 10.24 0.46 11.58 270.08 ;
    RECT 8.69 0.46 10.03 270.08 ;
    RECT 7.98 0.46 8.48 270.08 ;
    RECT 7.14 0.46 7.77 270.08 ;
    RECT 6.3 0.46 6.93 270.08 ;
    RECT 5.59 0.46 6.09 270.08 ;
    RECT 4.04 0.46 5.38 270.08 ;
    RECT 2.49 0.46 3.83 270.08 ;
    RECT 1.78 0.46 2.28 270.08 ;
    RECT 0.94 0.46 1.57 270.08 ;
    RECT 0.59 0.46 0.73 270.08 ;
    RECT 0.0 0.46 0.38 270.08 ;
    LAYER OVERLAP ;
    RECT 0.0 0.0 577.18 270.08 ;
    END
  END sram_dp_hde

END LIBRARY

